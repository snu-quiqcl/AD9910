`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LzK5yl5vGFn4usIyariozbxSIKs+MqOwLOz+NrjzoyeqroBM0xp0VSCNfUR6T1zh+lItOicThiLP
pYW03UVFyQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dN30TDCWlL83eZBjjW+7Ct0buL3q05m15QHd3KHRgyO9XPH3JmxKHh0zKQ+GVx2YfFfZKrXyvSw8
C0f/yWzWpB6DDMOfQWVyhF+GfkUaDGTtrIWhElNbq1nJR3thD2myK0TCHfwPVHVxzOGNY/8Ert2U
PmD1Rd1tcnOvMaDdbf8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JOs/eJ8nM+hzqsP4JZvqWCCZIUtoqXv1bDeul8F/o/kW1eI2ofq7sKP6TriKzJ2oXNsJBfdyrbZU
QW0aEp6IKIDmG5PwyU0IQYsFRfdy9AbwLpAhd9r5+3lXQeUytI/mMqhiWsR69FSX7wso0dPVaa5G
DqlW8mCikCpU0gAOZJ0lSRu60/PFXQtkF391kuuKfzcTY2tQH46pXtfP8phL7TxrX6iHnR4dSbOC
N2La6Jn+8zhjIns6txJCjSVp46FkhZIYFFl6Ywg93S2l84AxfRN0Q9s2fc7qCuB3Zr/C72/yFGmS
qjBylW97jBo3dF/HFturE82v5qJ6PUIAKZtsTg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o3MPhhNaSLxX8FcxwrYNVMwJJfdYGv3x9Jo84FasFAsEw/YnBa6RyN8Ep/Vi6YkZLwICX/jvVLqx
r/8NAPly5OCQnw8ifi4azQSNbRe8gSNEkPqlw6cqQUnOZJNDmq+CfAZXZtHfVAmj9mt0adCNoapE
zuckri8xnJRxzAve/yww9tlOOuDEE8DipECM5/5KAyT1nhM4estRoKTqNKsuqxUUG6FTWeyCF51s
FUCMby5+xM573i7RXGqEpF5OMLCUhb5HmxRJS+Cg6uyqrc/tGedVczA5TXgowGL7Kde8bRSqD7TR
Qqg6G8kpDi1St6Xzm+WtcVFHf9sZUZZ3uBT/VA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vBIzpg4CIC3z90ojxOBd+UnN/hwX35ZazMv4QfBpE21UYBVLNcLQe30yrAfxF9MKJIZGnHzyPZwL
g+FTYrLok1p3ojeUOOlJTEDQVsHAXdEb1hxpIkdVRTQrLqDWT8anUSg1DqWzBv3RNBDIMsBNMgbH
+bwFDwi8N/AYJAk8LQq3Ce0ffll0KgH/E07qYlkX2ANpHOzBTEZCTIIwffTGyVPhofaY+dq2SJGp
J9TUHzxJrlCf9veo8M1HnT25q3GYr8JdD+6jRE02aFFKxKm5at0ipqRKioEpWmxQHHGIH3bdWre0
r5gsJV8NNVueZLTw4i7nEPzyZ0nArjzy9LIIDA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qULPEY//q4KMMXq2x4Ww/h1G2GYGSS48hFt5qpfySwzHMslm8gkID/J8+J5yhNGfOF99RDW9ryHs
aJXNAHKi7IZleoDa94nTPLuQ57ALiajYb4M4NIqvZ4J3WDuKfLoNr+S4S9u4L0yOiwWIyGFPUQAT
KpbbhDyEj2023mFdlMA=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m7P2mzWmTOEbEFwkOD0Y2duZnShSBJwdR3fOCcTihVq0Ujfmw2VVYZgesOzXTQi498JsUYa/Qbx/
iUCpsPzfll+cY7RIxFk08xSFiPABl9E38UHtzD/n8vU63N4OTfWsIFFK+aocU7SCX7/a6yakK80b
3I1zaMuUTEFsmlXKGB2GMwq1Ixtk2C6aLg5lgj5A/naoTs6j/tnS9z6vn+htuG44TeDdRlE6QARl
0ig+WGsspWRyh06aOs9j5dIVqLwX/FPaqOYARnaEIhIAEarTRpZ8t4SPGmaQMKO3jQLnlzCrffrB
okDUdzJtJ+cv6b/THQo4JiKXI4ZBmwxr9amEwg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296032)
`protect data_block
TeAi/urTOSMW7Yj6k5jN9FzB8VGhI9dZvSBnTRgzo2a9vkD+8YuMn05Iq8m43ATLuY07/uQyhsUZ
3GaFgCGehOAFXlFk1lRMD2baqpP11O8RrUWrEg99JVVuPTeTp1LRKl7czP84JAERCzQdPWFTy/xz
dlVZmSj4TYxgPYm0ERrVRDTzx42YxRqOyXE6vzCMxMcdYszWyqxqp1r/zBqFbp68G25g1UQZh8gQ
PzeSP4hJxiJWCZb71CHmPh7VOzYGfxBz1X+PGG+xs0T0KOwlOs9GmNRQIdiCpyq7KLqbnkDdVCuJ
FBedPIkyNzDSqCZ0kdd2TCkUYjnJA3Q6dNQxTW6PhTsdYZKnsvr3x1qYELOsq+OKDzkrd/gqPF6F
cxiV6sZNzzGK4qvKgHtx/HvyKXvPJPAqUM/uz7opQKDJMENHcc8/CC+3wBiHcUpgDT5YVNP5jtY7
yK5YwbZDVCWpNU8uOyR7qeO2+M/LeusB5nbMczBRVGhVjHg2Erg4iGYvqhWtvC/IEXZDOfN6akj0
woYpTKl2l6U4M3WpNQkU/+nKmh/1wHmIOmCdgnL5FjwcSZQuv9wmlk4Han5rWu8mYhYE0Nog03PT
yz+SMD5WmqWG+izhp2W4RCIef8BJdtfmrpH/gE6paCmKsiedazQjI8JD7OPG3ewQmVr6HszeTZDl
J9/1NlDu928DlvbPSUH/ECHR7K9HCw6mXCOLE8AGTFvagnxgLqQzurmWNaQ3DyYL8J8pWK1ftfLX
N4y7K1BF2Cgu0j76+2ww43gJkY55y6pJatRFM3gnsbk7ph8af5h1h7PXeW7KX15uh+ozEa4kLkdy
vwGB8I1ihpbS0k9lCEELnB06aKdlkhsjsiggY9K6eDFD6LSq1LxMpa96mOrHBqirgNvHJqcZ0RnJ
1/f1TXVrGVXHfbAdEmtW9PNqLWfaEUo0B3YEky0al9tUveJZIY9Cv6zlRf/NEzEwWFYRMHuNgwl1
rH/PnrWpdghX1N+ZuSwFwywgtkyl37eRdb/DKolR/yOhRNrO0zxTtB9+lvzRffibrKw/JKPX9R02
hppvuVRf7rFuWGQgCIszoN8h4jwBN7U9aEwSghIGTPJGqYP7z+kjK0bqeD4BJCPKESVpuaNEssOF
9pS14bIEBXykl8f9qsfdew+cxuGgbEDJFVgUSrfV98FJmUVhvuSETMoIvrYAei2eqYTPVO0PSwE9
N8ruhooPz+eomyGqNRMD3AN3lAt+6trqo58uJPEjnxBzAdNYO7fdOsX2J4qIvnDa0t4Q4QAciF6j
MFfrQ6Z6VjDCFQMBL3yU+y76qEtv6PiJ+KOg9ChX4WanF9AYy9sb1VO7rd+09SP7f43gYuB49SLa
7v+rT117Q1L4cWv8McKnzc0RLdi4Qlh5Kn92HvcbZtGBOdowbrxNb4CXFnhNnFkRMSxJfAI/f87+
/403SOVorMwA9r55X4ghW8mB9vvuBhrfC4ZxI96+S4Qj02soNwoef1+aVBmrI0x/by8dGJlqwOWG
UwQqySX39DQ0mChrTAsAwLU2KOK/f9c3QL+aQl/DQskN+macXnPpiwAXywUsN4i4dxddjo8RiKis
k8pAWfTGoHSBp/is7+kMfEedZYQbdpuOvf9lD9A8cmppFGEQC4pzyDZbfhfJ0da1OZHqR55hu0nS
7H+7bp17xQy6t7HIw1sNUBQRQmlnJO82onZgwHFR7Ufsmwd97/Id+q3yMilkWT6d6FQOhnBaJzfn
3idAfHB1mD7jZUMIuvEuUlyOwgcRRPtiuAcv4/956v1pLaFJqF2f9v/3eHrglkrqjc3XQIKAH+Dt
9XP6mC1jAjMf8yMqdbWDcIG2qly8EUNy/HizCnGc3L8iGXTy4IDvQ4rCxlHwqOEX5BesRo4yVbrU
XxWH9XMcHOHOaYU7mjMlwphCu5IBDAXCwK+kzpolZb7JMd/YxP9fHeGj4m3cBTJy1RhaAZY3ViNJ
mBqnVyi2u7jfcfw4gjAPetiEMk0m8KyWdjzbPbJZ/legJVxb9wPmmyhc9sPXgd67mxDOENjzl7mW
8ZKH/Ha29uU9QT4jfQGP6dZwBCeweQ5GX51K5kIXWyNzk7L2Ahz4b3TByNdzN+biqQrBb4eXMPpd
x7hVkcdB+InPrrMh0TXOKjoDU2AfzHfIcaY6oVKG7uJqyM+atiDGpDzRhgBskWl1X0DBgGS8T8g+
c7e/lUT6OF3uVB1PWzryMpOXLhZub9OUSxUDuCYA0A3PE3WL5/E3xf8+Eh94nJekOMC2l80wGoRy
oECGk3o4eQtZtJRioe1NmxvdwZUu35wHGWQLStoEdHCFZf133rUhFYcXqYlmhnUkUJxpDAU166xm
WQrpw4kUY5JVFUwkhOmo2ivsJHv6XrvLE1dex2OowIx2ns3EO/+Yev98kYRuGT0vX6Q16JKP2NGl
cQyLCjgC++Fc8EW3nUU+UAjSCjQOTrRH+aTRYoa0sXDSX983egSoTVuT77xLPHFZ/cue2z9oYtWI
l2tlR6NccUivepTVhmOKa0rKFypSzk9+WmD4SqjDtjZGQb6i69J7xcH2L9mrVSLZm7IWzcMdCGjY
gkQjREjXZQMoCQkZ50c6UzSYJTTnRkc2uT70N8tw2noH3C9KR4j0RkagvuXG1MXxFOXQupT7bJQb
yUm9Q2un1jX2GBlewgFwByI0tKWHLH4Z0VzK5OfzQdHxtWyGhBIHsfFF4Aw4qmxKqYL21hBsNxUD
ng9ncSN5rM4pXwq25nwIQU8v+T/t2R9cStoLtRLZjYe2FTp+ljEMUCuSQ86zyNP6HmbYH8WP6Ce+
o9ete6FPlLs7nwxSoHKB2z59LcQ1B/AIjkwb9ge9ei41kTg1UduP3+POR09ylpph5+zl66C7F60I
wnN+CH/dWH6qL+C+rwlmteMZoJRaYcOHb7bZyfzDKB5L7WgfBVaXkUTLInIBGFZ3UabHtwI83hti
xQokdjjrMfr4ZCMafYbn9Zvs8uRlMbyoAwEW6H68crtli/ZOt3nU+2KGuBhdtZktXwx5ImIRDYwP
g8akn+yI2wU0jMZqmJsbNlbxUuWdQQDmmbFBLaEs3yN3wu7yP6iy4+5Ffs/J/wFnjffOXOU9fhJk
YGAyO8J35UK5muaxeI61r4bdKrL8G2PQgngnvsr2iood5aaL+idp6vkrWWxGQ2x5aP3gQnonbspB
KHkA3Y0IHls/QoHR4tGqlsKtQIAMw8XXthTcdIOwhVKsuQIF3DxBiB/h7faeJinU2Rzax6ZOLPka
YgMfy7EP+z2tMSLIoXyGjNBMAUhvTJL8llM0gVuEmkDO1ezUHKAIeTdMhFcNc/cnx0Kp/D1MJtXt
Kbhf+NI7yIpS/5EqMmOCkzn8Ga/J+xLimGQJ41OX2F0EPmxb9inzRKh36aBZSAP9ko/OiMqjOLIV
njQxXGcITpMImzl++5Z5h6qeY5w36TDBz0+4vxEAJnQGHv8d56qYAXKKHer4ZZL/fi97FJN+NqBj
4ZxlH/WBu7XcQJtpxrDFRX6m0LaT0oQz1RPdE33XpR60fcp3TiWwgZUanjn5mna4BopdiRsalZnn
Lj2faEIdQy57GkSNejJjZSPvK16YT3wvXyaUgbN9MU3Oe4YV5cDUKDVuAIp1gSsf5ai8bPkBjB9I
UXoZYELlgRjzVKde6PVbVUICmZOupkl6dd+uXaf2KspJuq86l5ToozOucpxdHXE2DoQVv0WSf3g1
saumPFZjweui0mgsSSpzE3CYP8l3aGzI3LSLvjKFeaVdW4Mg6Ld4S7vQF7/5kxb283aUafPC8o6N
aZtBDQ4d+V3o+rkiUovWFcSk/XG8lHf+qoSlEH9yCuEzWcx9zJquIk5B5hbmAiJB/m7E3M1nL3hq
pa32IbiWfRrbFg+f/to8HCHn2YwAUH+caPRs4gnK7IX56HyviusODvSACtoU3p17xLNUwPpDv0ri
eMb2DHcr9tfMFTo2dn9UIKd84uq/S7WspiMTaDOAcohE6WqqMcXcATMkew0cIoL1ZciG9oM2basA
bs1vT7ViKLZg6XnuVQVoR8A9cuF9oV+KsZSa7ykb7UtzsPIa6IRcCB/TaIgonbUZUXLdfs9MbqHU
Dv9KZvqCWFi5uXbIq7JcxGbhN2RfhdnQYNrTdZX5uQmvhFvAFoImZ8A/uq62+Q7Te6ibsjjc1gEA
/nbdBlwio0h5iZ4FFQ+59OKrNhsARTW45PgK/zOjUqxiEUwIPGU8ELLhufSt6VnIgoZkJBV9XXiE
wNfGHD4HBvMn8y7OTKKAf3D+fbf1+tZdXAj16USHUlF42xdy35cRD8mKF7zFeyDpNeRdCJOLONGD
Lq7MjlU/P5i+u14K3/XGQaxJymCGPWyiIwo80cJA9gnPE3utgBN5m88mQyD53TcECpkVZqaetwY0
C2VuM8Pmh7VgBDtJHt7hXUALIQLRk9uHO1is3ZRP4aHflzwmaGWjajptl9Tju1XEO+fFpD9kvJGY
P9BXgVTBAtHnPSm8iKSubAVa8uf1ujv9zXooWhTwv6TICzhfpeY6gI1BuCDbDEOYPq7VYkyo8cLt
avqmxb1UVVRLA2cObEo8WE0qVH1x+vemTaLYF+MYB1e06zpKuSDczC7p8odRMy+58Gdfu3KAdc/M
L0I79P/32LAduIsQyjc9mK/utGjw+rmL8YflDY1wyTrZWoStkl0WTB97xPSYCslx8oFPySUfAcfg
99bHKhlzRN0RGhYV+YkqopOikt6ZmJbmf4wGha4zbM8QtxSAuBiMgFN5HbRTqLAL/l74f5L9n/jA
goZ9/AwrBVabs2O4bl35HAJ8hTKjbVbOUE5EKk2gq064gMYt+Q9XN/ysjCrf/9eUkq6Dcd44GX8e
BTd2zyla5A2wWbs0KtWjh3cW8fhychaBdReVXUrLlTjoLAGAdXWVm72DrRx9rzGhNbpybR+NP7Pk
K0HK4ErEGG7TCcInKaVGoEX6IvAjzPwX7awJXgC6+z13Ec+AJt1xbFx4LxsEvSzt6xoPJB/lkj5t
GdhhoyyQFu0pMCgCNzLHnHvLYllQGigfKP2iTnsWW869gJ5HYQXlizotYvsrwNTpHY02tK4VhRGm
KPbWrasKoIyO96dhxdw/mZos9l8c+oEQMynrfQEVrVml+xuaVxhtwR2vSd/0QfX1fQoSLSQlpFVu
MBqhjNsQs4822cU1a2e5+PkD8BFZHH2AVCX/lBD2Yf1eKz9QeYe2kWr5iAOaiDMI06z9LcjD4LdC
byJKozi258+p2fZSu81AU5T2fDwjfzFy8nGOjU5VY3TNVCC+WrP6/8A4mJJ1Cc+YOEfTg65ZTx+u
9iAxdfcZJFwB1rh9Qp2kWpv3+lqa0ZoLN/B/ZrOcoY6dHyApI+4SUB3cU6wtJjonrGF5SmUw+Zoe
xbrbThMMkPMyh+5oK8JIFTB8ZutYt/hGrin3gKG9FWys4OgAHUSgoTIJBtPeAJ/L9/l4W9zcfM74
uYS2i5iMSuf9a6eywBakyUvUTli2zTu+betQH4eQCoTx7gVzu6/dpffQNRoVUp+DqDiZ1dMLLZ0b
UV4EXG8EzWvEVe49hpAf7PgjGgIIYNznbKgUazCjH89XfJ6WTTmmOuVrHGIM4pRFE65SJqlTwKpF
1d2ej7raAE+4AikqP8UKEqImXoNX8MkiTBw6Qj+ANM3axAjmDpZhHAtoVF7HPwes4ki+IoSGCWZ1
SoBWtVO9T/DrLOFKo8sCl2ltulguZ+Yl6PNNeTleTvFed3ZxEKwFoQlGHHFlgo7/ls0CpPvLKUMY
vWB7g500LRqlSQeXzvgUi7P+pVdpP1YLd27EpoM64m7KZkOokatqoJGxN0Xwlzd4MseA+OO+11O4
qhGnBBP24Tvb+1eFW/PDNz7hl7EytsOu0PZ24DVq7mIff3Oj2SefIyosOHSgQGkmXj3jLCKGGvMy
WwSB+jDobohURp2a8IyJQXwIdljAbbX6ipqNdjUPOllT8Xyc9GFeFr+ujweL5IuODqnaLvH3VMEG
7y5v5338bWtTA+1Ga+EHXFSsOuY8ICbH3JDQPZNQAnEKg6gl5N/dGpfp0pHuquBymaAg0jqC+mqA
s2FvMe1ZLn7zeJstfwHEshhVcjOyzLTK5jEjrOtxx28SLOlxtSaMi7mZc+JKO0sD1AN/dSQeBP9n
/zue/2uvJEGJ+hS/ATllPsI+s8j1Uz+P2oVAFgGF9A35ceWDpTnkv+5zuZ1B/ODj7wB16Q3uhZnI
Z8Ts6Nb3WKMEgcVps+lqtgHJPI+NE9n/biQVJWATVue5CZCiM/NlRcBSd8sSdikRqlMA3Agu5x8z
BozxXgY/LON9ZFqJPR6wow2UbnHzBqrlPtElevHzAOlp0ivzSACsLfaAkvOxVyYunO1xg3MVeuZg
hxSamRxVaOTyC1NyCZO/VEIMdDWPcifi/Kom0piAY59IAVSWTec1xPMJFr0+O3Qc4UkDv9rb80X0
B0UAl5whVl0QR2OyjPjVYrCVtZr9qF2if92kG/RAyUpPOAwGlhmRnVMLLE/LtEYtM229/gSjccnm
2t7uj3qFXh2bZKMFbXLGJ7MkwBj15gMZYp+fe1m2my55x3lJmcYs+fKXjywlYirjAN9jjNwkA211
YJC1oOrofCFsX6oNBajboXDVxrIeC+Yo3BVZeTmboXfQDBy5EyzzL97fBiWxhLkpw8oqYXL3uOFA
9IPPV2Phkw4et2h1B5bPz7Tzdeukd7oxNPglfB3IkBxQsN4JTRHcS5l4lpZ2aTM6Rerx55WkFt+j
Gul3z9OLhRVdI593SYLy74Vl47CBr1Krui+6CFa6BHLSJOZGlyHPjYp5/rPFrQMQxE0JHO+XRb6p
PJm4EE86DO2fYIZMtvuWHa6kTNsjAPpuJWYMOYc1rL/wgBeY196L2jQ9+M9wU6MnlcdZNeyHWo+3
+T9jxPi1iEZNZ3TWmttpXQJtXeEBOvTuVBcNDp0eyoZVtWkpzGk7xdCWozpxoZ9KElpt9A6hBTU1
shKCLNBHnbg8oVOFM3aMhgYf4Iwxjt0rpXRdWcW17OgEzOX576klzY+6uL94tQZxCpFWkisSAzx+
f4iAvTDVSzpa0kMHju3IuDG0lVC1cZQ8T8QT9znxGsCJLkesV3dzXGKXAJvN2fRSb6Vcu20f6YQ7
DoNQS/qmgG85S/4PDA9EzcZb6MEpH0ESFbC9wrFBDbhAPE5YlnHm7JDDsXwQSuXkw0II9GglDujk
he1+Csdc26cC+dUv1zpHumVEwAXwzIZvWCbydDtFDbX5Spr2mK6IADWTUzY4GQPTIpkjTOTJvkcH
zrMyYpWq5qq+8sLMuhiJziDLCe4XYXe0JEPyMkl2Of2W9XNBUaKmFaOcgzjZf/G2l9mR4Oth2Oyp
Nt5hBw5+pprHEmRJaUh9ooj2AzSzDmg44jvDOB7G5smDNdU+uGx+MM2gzQ7v/U8qbJZNYPjyZUli
gN6hMaozpQ5ZrWBco3gd1lrHUGQ7Bu62IWiEEEBE6G29V/FhVrAX5LyKwfVOlFAdFhq1ll7UMW47
KbHZ91DY40/59OgdxFnr3Hqmy1zcQ+WvyY9BMXOeVgqyI6NrO+5wo+d7jDCziStooGEM1bRBZUrn
iPPoaL4CgDsO3URJ7atKjC3tTod3+bJ+URZtMliL90w1nTYvWcoDAPDDOqJ7Opx+3nOq+xnMAVNH
mqjoTKNpmKTEU4wxVlHDM5P+6rMqLeIrSABT4YVULZLwqE0c9QbXrTMgDxdRBFZ/QgQtpAjzjpW3
0oix5SuQ4FVx8QZLx9DqRWArq2iw5fh/lz0GprAXSYwTqNR/XKvyr7CJ7zM3ZAs5vbJ2NRD6fNLJ
FmXg1Uj1WqPCRzbAMsmd6svkBn61IKId71dEaQOf2KdSTGjqyic5a0PjH8TIc5mcO9N6gDWy1vab
UnMTjI8+tnIdfqDKtt02OpuRNl4vVjjciI1PCHPMwh+hVvRoGi+r1XyMP52ACUwC/vrXFTSLu0VP
vT8N5Uzi5qUE1nrhtpvG/PQ35uFStWcIAzRAuF1C/tpq30Uv3ZuAVzrrNbhHvANXpVQsUQ+frBEt
qCxVhfSPYsadYa8GUlG2+6YJ1vXqF/lik3blRoeOmbMjzogTGAenZ8d2gj943mpbnTMR8ObhD4lU
xtuRXdrgXKlRdILW5lRYXMvcTrlFzTrEwon1WHUZ32EZy/qJ7vVKtVfUb45PrkAQxn8DxeypfFz6
Gp+WKgQzbsY0DjJhBMoIMEQVq52iiMtrn7neOAlDgMenFin333r1MdI/dwsC1/LFYI+KwCedKAXC
i/+ETY/fcJP1Wp720q1ccoJ+xgiDnwSwEQ6ri3CuJle7kok6ZJxTTwqA3USfw6fTwfTDTXESVl6G
NCfMnDY417FIQAABXQGUvN0opAhWQ9CNNf7bF2dCDzekMPUHR22jP4EfJ8ozkj0qaJ8YibqZPqVI
b4pY7i5w9NqRxx25DCyNy+h1q3bIJTLer2pALWocHGxGyEMqh9Ks6oJfo2pFd8Kgz9ZaHsbCSoj+
KQsNvVDI3N+G8qzrCdt2n9jpdnM4brUlubhaiMYvoww3i7oPbckT3dAmaPXCEI9VS9kDW9IgiUdf
HgQiXc2CaQCVlWQGhIDtIslLzEbDKl0/NEo88EABI8w1RzuK4sZHoUY8VGxIgDLFGUfa+7luvoTN
meAppVksSkOOEjBaajTlVI4X11AwhxEZthr5e9h+SeAJAUWf9/7OP4CooKq6LUzZQr7B57wEpkwv
LpHX2R0MytamG8gu2TwBBkujG0C+k/RfNDQn2cTOth/UORFnzTaXqwhx4k7l2UIYiuJV1iKTWE2f
vlWubt1L2OjyPobGpdwwVRZJGMEJsM4cZ/X0F3vYez4ljSjy+kwXptnUt1xTydh8zsJWEOwjRW3E
vlwpBpUxQEDs+qQym2OQz/zaolWzouFlbFHyJuo60hbv96XJV7hXc9zXgsXkhDarob+mg7D/yWX9
caTSA+2DI7hyOWAPJjmY1rWZWnTY2nV328FlwsfwT7CjvVzC+3mHpGp+HLJkEcyvtz5h+IfXZ0mC
/2IOzJRgCp5UPxIHVlJ5tvTdNO92rKZ3eCExa5fXWNKaLO2afolqdt8WkKxEknDKqcH40HVGp7EK
45XP/PxWuuXPqzRVYlSV+vhmyFLwBCX3o6o9kWTWVLCyYH9dCRjI2W/M9wYBJI0AXgXnW03Impmw
4qpJmI/8U0/p3Mf2oyeDEd0rIP7lvJbxdqcO9Y0i3aslef7QJYG7HkgNbnQNscrndH1HrsZqap1A
VTUgIp6ZybgJZtyQkuYLEv9MWD9ZzsvTVOiEhFAf2rJyWYgFjEyQv0O+dtqLr0GHLTvSiEJ8DB8I
qc57L59psSPhlGa8iP/JjLqIBWD/hJzMCl1qDJTreLVR3omu+lxDj4AvvLcpHs+VMN1hT+hr6HB4
cadI4Kd2M02fT2+6epSSA18uJlzsMmiL1haowEYV5MzEJRObSS/uFP4/IBkBLPftx5y0gK/Rjw90
mSQLfhdqlt5TX/OC7lE9GhL/LsYgBF4S8mFEVu5ZtiOJRhJzN4dUW49HONjZ61PglZt7x5XT0jLF
XlFYfC8daShJSnpqiwx9Fsin1VFcYHT4jNf+ZhbxgN/PJ2UtPe2xHPS+eJz/02CiZLCtgBMC1cK5
XnlDHNTLXbMZLHaSfx53h7tmWtbtXoDOru5e9lI07HlJSFPNzB2GfWhYmsQRUXYOCg77gIMMG1h6
bfC2ClJf7Hz3iNzZkPeY06ZTl83N32f0OOAplUH3uLraeFzDogVlgDeZs0wOdQRjiEhboS5vua6T
TSTzK9BEhk8f0QoY7rHuJTg0k35F02avHxW5EgeqXSYiETRQ5nwL6A2DZ7G08GA/m3etVDxNCrMB
WLigSA+YylWkyUKYijG0XqgtDFK/jOHponS5GQT09S3B7gaICnRZBGDFzj13i0LaqEsi5Ggfm/pg
VdlKr4bpckhEUWHJ4/XymrHqeWJ0aP9ZreslMU5utq1GVvUnWtb9IdC3hjNo9g41mZzvO6/e3SWw
v4JwEMFmnyIAztByGyoBYSS9vGZ9PUVM6Xd1fBfAsqez1p9sUoex8D5Dg5F90sNhX6YrtT1kUOfV
92DeDg1Enw9ZjHg251+cyBNvQgfhY0CST5pjtqQxn2OdJ8JEvMToMYRS8UnEpNg4q8sgbGCOy4dk
KRq6o6Q75UwusxnyEsxNV5CtymWrcXphla2sM76L98qJ5AStSswAhdIikOXozNi1fYiu36dWr2Eu
K6BHDswvlybKG7KoSCX5zJGWG/cNnc0m0ltklLzEwJLxONRHtCq+ZN3MoiHSdTURfajL4XUWL/mV
d6ugemgNKi2yAdwlTeqrJZmsMDfypjA3h5IOFeEBe3Dj8ZPP51Gc8NSkq6wcoJx0ZH7pRxBJS9AO
LSBHmEgA8ayKz7cyRyMWpCxkbScWX/9d0c318TkljBZJkkDePu6FEqMY3iv9ZPO5Ag4p3+jiKDwf
7myEMgXjY6zq7XBQf1ZcT0UPTdpZ7FBjlAYAepyjOQSyhbC7lH6wtvq6HC9HTlrroSd9ggQIuLr7
X9lpP1RH6lpWQ1QL4NCz0z84CPcA3PWVUMTz7tpMnS1Yfst2GBK8KwfTXdvGdc2dje7HAEinM9ep
WZujjfnZS9FMpP0iIsyIBpbmy4wWIL3P2ATaFGVy7kUlF2xOVRtAWxQ6P9wlZoq3rJHNeQEK52RC
P74zY1ET6nl+23vN/YkOyNGTrJzZQuxT0YCdCBRmHa2Od4/FUb6fFv4D5r2wwfx33VmTceQrwy6e
dPH6FzHGRu+Fv8LbHCb+lJS2utdaVmOq7+xrVHVyY5giI2Xj/DyiEmCgvx56ChhoHmN0pqmUOC29
Auqo1072yU3KevfXhllHzm9KDHI0xlqraN6wcjKnSPfbOe38ZGh9o0yegwHNyXaFNSBYZJzLg51H
PWwWaOJPEkO0+L5igYad3esrruotxKJuMmdIjLRqahtfo5rqcC2lbervjLHNMmsdZCaDcSv2tPky
E8/EUsjtUEYXsvVlhBDYVT1DQ/UGCHr5Cz2JGTVnF3EmHte2ryh/yIsg8xaCC6O5Ak4x2urIK2jy
bPXPBO/7yZDZo0LJHpAhuijRKyGKLIIjdBrLv+prq7SpPw/6aX/XCjiUBTDfC5IREBl6uH5GceTi
xx77GBFb3fGyy1OPG3jtcokRcjbbXZGJta1jpIG4v8e5opEhPSvGu5+fym12w3Q4dRrQuk2H9ilj
KBlyJ061mAHLJ9F8fiEYKc4+4zIMEV22CpKuLbxP6GZL791EeK706EOiTe3alTOz7n6Y4z1KikWi
Rzue6YBT/Yj4VYqWXF+nXGK/n3BLa8vjH+r8KuRPzrcBooJhpD4581BOI1isuZYkfs+n7OcDlsPa
U1RLMWw6i2AIJH/K10w19KCY/6jMhmJRVINIIfjtWszvyuJ0JGLn3bubdD0iis/4yh+cR47ddPXE
uxAGPGYCuSvpStzmJ89itd2UIkwugO4y02Z0QKZU6gAnIuU1qYkWZqCaSpJ+yhgNKeYVvISvrutT
rm0UjT+hY7SNvmaS9vlSMcI9LJRtM7zCyHzT6lryiysT2xzAnX+eL8Sf2jwjr/FrdlVsWnUxiDST
AizSWtNHfnYkp1hIXlbcAVQA8+utiACAr4sQ6dDcC8L8WR69LiKXU48nqlZUqFnmMlaTvM2rNkEd
8Q0GxOoYNtPI81Qr+XOErVfasr8KA0kZvggcIKtTk0p4aHi/+QEtFudVVeouapuEQXKk+nyb1pek
ed/NzNOAQlUizzbdbBl/+k34lfGwFypafN852n2mXCLHA1sCHboWaIf4zWkbbPwVEwv0MHO+eqz9
8Tim+hyJ5zKoe64xUwEvo2PWMuUwT3VvhS2GYoOsJ3QS2xPFQ0MX8vWwjuqJ+u1cu9Ugw/eRd35T
/EEfS3iIZ4suZzSDZ5gzLEGhRE5G7s+oUD2vBCGCVGlrL5QsvIGpjnFfIMDsqn7jUjca9atVkSjx
ft68HHXdfi107j2mkC7m2Oz0sCG7UPo9pHGvxQ375E9cQU0wSvMVsqEmxQT92njmYZBMk7UB7tpY
fc718G83K967KPPlH2G/g5wUMqH6bNUgEERwka7kaca/bQaYwgmFwpNcL4op8wbOlH1pjUObkdkg
FW3IWAx/DfMfQ2VkjtYhreJPLhha3HylN9xHVxuEuZgavx+G6I4ClPTBoxpMfX0SKglOb7lx9q7D
mjjnEjGavClsWr835kSrBwAsSfe7SAPudOlqEV4VMmHU3JijV5sA2uUYVqz3pAY8C7CqSIHcqNOS
hqel64vXRDBO/qMo6RPSFnDa90+VfAO8ZlI71wBoku/JQ11Qh9c52g4TwUzvXOLgD/gq/pJm7SZD
qVwara1lThfyoaj7QRwqdbsKk60CdwhBKFRdPzh9d+3MqgA/iH0w04FSh4NXZToH8d7xUHUgUlxK
nCvAtLixrO2n9rWbuqzbEoMTK0uqO1Racxv8O554wqEumV6PSoa6rdyvYYUz52cEUNr3D/2mNk3w
U8IGy9gJe7GnppaCrpX24LN1pKO5k7faU/XVwzxU7WO/YotA96O4cXrulAsg/S8BZzIcosn1sUQ4
n/DpOFNvE4dFBvIJ8YsibYa5dBVO+wc56uydsL54xesDnXMT59s74yVBFJVaxsngiP3Uo8CQwIb7
BHdh7XT29SA42tGZ1y5KfzkWvlcRCry78BwZuMWgYdmfD98FniBww5smf6h4trsov3Gi9L7NPgPP
LEt1rpJBjLbNp2ECYDo/5HsKkw4CzzHf93fy2TJELTwNqLgOWPEAXlC/yHMkMt8F9MhYGblxpcSU
xWb/7KNUOGQ9jO+ghvzzbG3o43mCfQKgngqIVW5I2LroMqGmDPeJyoi5hjZNx2H8WdoZ8ZUANBlU
sMPyvfeZvrkb/xXqo9LhDCdD5tD1YDRO1axvU2PLy/pmywOOfHz4t4snd1I8MkD8Mh7lzzc73Jc1
nadTt6Wnz2FbSZYEyRjtm5RrOd99Qb+9JLiDcDqrl9ZzeP9xcY7kTbWAIph/qNT9lRZ/WtCvno4H
+kdjqiYYRRdO+mk1LYCbBNVhuWwKN2PIQ7jnGuBBJlqwu4mkFJk5krOFWio0f9fejupcmn2ZQoPo
xNftOXsKLtvv1JUh+xouRhaZD8ySNXQyeb4JDRgJwwuVadVwW95vPDHDLlDIDSQ9d2gu1ydfuzuo
cgPwjLWywU8znFO5OTWjghTWAJflL1vAScufvwTGlOcP2WwOa6UfUU9XKdbMYYNMHLA33IcUguSr
DLHhcdVpBqO2sagnqV8k4P50LwzMbeoDOG4SF2S2OSDNrun6um1ffh/pgxPBY2HqlEJTqUS97kJT
P/GNcvskEVO5DJmaKGRqxyTJHvpSYlwRZTCFmYJZoRIJipGtrsWGOh4ixwWl/fWE/3rlDcWXkElI
Xz0R0K0v/LUiBN+SGjkNNb39nztab+mri2Oll0iNnOY7Jz6gk6ymOvbgAmQ3W4z7kmOZwHmTozmg
bBjyhz68EFi7ojqu2BAY6O4gr//rgyRs3lxwPhBXmboUvD8ZDZsLZ+F7LgaV642Lg9QzJu5RqU4A
b5YLw237SxbF6GiysjVPppoYMAu993BlejhcshrUJNuKT95rC6yI6tmHqLQkulr57qAszPF6WzUV
tddq8QtLeT36c+WVuFousgtfwgeHmyj7IIvtbZ7PuRVcrDTJ/fxPZ+XVW8+ICfl+/rd66PEoyiHX
Jae1M5I+Exvz8z+9o+4a9Fc8NJ4I8UGNZliJfcj77Oita3yoIa1ZTQOIWHjQ1Hw9CPoE/whC2P7W
Kcb3tmdamn14M+kR3NQiyUE6ZslEOD+CeTI8XmsD64PeEj3TppjlSsARU8gVCcsN6+do0bmtLcFC
cVaSnnhE+ULYiA+9/8sTXSaHF7qiUEGCuUQI8ey+CokrKfnU8XK0KVxkD+qLolYYbbyP5u0Z/rSJ
hJUNEfEP2kOhW5fTOH7r3MSES2dVx/eVxTjEHM0jVLiwqflevNdU5ytV+SPOBeUiqgE5KxPNB8DQ
Wh0Mgzs1oW3+N16gzQ86l9zeYKOHgj0oND1YdQP2mtdvwJAjdlvXAoMXqfMWbQCy7LqKePFptGTI
l26Tl/oswNwKZbj4fFaq80TFjP/dxx0qns+4az5ajU4a3PV0bvtNl6JQopJsae22ROhaHInpJXP7
IPpWDuiBd73K0tBU6voDz2ek/3IkYh9xSH8ZcosU3EmB/oI44AIXJCBl8p5NnE0/99iTByRTy54a
3HwJH0jItakgqAPvsJTxBRxKeIl5yRppmz4X7jnOf+41TLvK0y2Gbcs7rIRi/mryxCf4WfZ3FOPS
WCaC9jr9w4U+VpaQ6ON3Gg3zOLMbnRMqxXooL1VkA/rLqRcbyfTREzVc4BkEsvN0SMS6QzzSJxMe
vgN7/nTK6giiNPyqZnFmiVnQ4Y4h0pcdWPBjrKx4o3keJNE0lvME/SA/gcKQRMUv5av3xnC3DbOo
ksv3lHypUGNYHpuzpaGA0pcrWAbrvLGZ6RA72lWA7juKPZbla+vNa0ZhWzmq/7Hbhm6WQ/GfvR+j
5FU273vUX/LI0GP/CDo2CZ4tITQWsZUfTdFOOXf1FrKm3Rnd/KZwQst8OQX/DIcSsrb/DlQScWZc
TFAyQPqUaCK9PS5EGfm1FnKbMrkLdTjt8Qk0B+E7WYJUBll+hNcKARjf6j+oLxxc8fk/HhrgJ9lv
kjc0WS2XCrfeBB3byHNPSbWgHMMlhj7px05emji1hDKOZvVbu/HYvHvVGvAEmVtcPdgvUVNX9ePL
ocOePSEHTfxHSko6KE7myvnA0Eg0/onY4xTI3fJuO/0oAPrMA39NVN0Cl6ip+XlrhTXA0T5kvHqS
NABRGg0UoG3Jh3JwvZDwTaBJF/Pmkg1rTrnGC8k2u28d5uwBd3UO9jRv7Y7IS2KNNoz2oTEpGFRY
U29T+C/4I4sPPnNx7pJ0GQeQc3ZVEC5lMr1pqpc61tYec6aF0NYbfQ/I3IQlh5irY5E2cvGG5IQH
IFc4zHjxoQNli6EIlA8lIYxGvsTdSuMGF65EEP8TIQfgZ1ZyIS4b5Tp6FI5WJj+DuCtciNqe9mPv
b0SIxvDk1buLj1tX/s6nRof8Z5p3n1fqCGqb1Jmg2OqynM+J9xHuqVRijZ+juTCHSmhoi35B75nZ
GRvkNraBIse0HPT4MeRiKOyi0FgQLGJIht+mGMNW6gwytiMJxsWb4fFi5EGNnyDiygXbVpfBx0Cc
SEOlSeQoNlMiCSBWlkHGYcTI3q6pErdesVGhrS7jX7einYYNcCxBMFDmdkCqh6wU/UksTHI98sZC
z/9cc0E4UeuygfGVfbyssNj6vNEBe7DAtjjyrdKxX8F8udr7IU85eLpIK6xPIkqos0UF+UzR5GLx
acEaoAlpGbrWbO4zvQOyd3JXkLQNyc3e5w/IFr8YoQb2GwBznQGvL46STVhO58AU+Gh63Y9nniMN
CppUa9TQpfeVvAoOY6FFybRLZJ4R1QLEMDytudxmb/3mUOhGj/LiGohplaCShUi8FIcbFTKAkntP
WcA5v1m4HVY4ZhFhrqObisyE4Q+9m9iI9swzkRyvO/PUbPrp6NnjZip/1NT7naY/5x/18i3GzrU0
21MCZhxd2g7SN6xsI9SjKV6I5Rrh1h+eX6m9bdxCyrXMUM5NHsKgda26VtiKOsp0i7HhLnHE1W/z
KtRyl2FZCfBGcvJYNdmmq+5uV4NoJwBPY+lCNp18ox6b2wgEcgABP7JB0Uon6i/PDecwO6SW2sz6
CAvN0fSwU92KOJfEpT38SdutIlonu/K5KSKvd483Iom7QBI6w3/gLZcGEN7uE4HO+BSZexL1sjWP
ujKR8Rn3LsQAVijEBpGqEpYYCteLF1oFD2f+SD592pIxkUa9XofZ+kMHnoOiTFRsXEDeRkoFqhZP
2IGxmobKqNtTU0OM1HWEzkr8HyZUOXwv+LnNxKw97iFh6Ug+UIzbv2xeEaHoV9VA/U7rvwNQP9nV
xBUtv8W1MyQXxlve9/69IEPisK5dOsoVHn4NJ1IEaefSa0k0rGgfJKnAVtxSFTJDsfEnSrLYHG9Y
JP179lADYCEtz4LMZa5yZwk39Ift93fM0frO38kK9xRvVVOvCBIESAfZSx9tTSsnr2oxg3qmsIls
75YY0eEfdzWJBruaSyht7g7QcMx9V3pcde6AFvc2OPzlw6Oy8yxYsOI0kAFfw1qItZnBAmJQCWKV
R9xZqEtiQlG+rexIpt1ljaYKOnwJeozyUbravOSeGHkF743KUkc/EqSEYiPmiD2m7GFnw4YXorPz
KQSNF9V7IuG9qiR0XrQFBmwA28A4HjDqGtCM5ovKx1Y6/SGpPXOPukYjbPbmv5g1LHVaRJ4Pmmw+
KVCOqYq6WlIK1+VQdPrisoH+xBO9UHoPCM2aDa50FwdCFBwmSi6Abq5OlmwchlAUfrYLMx/bvL4x
A2lmQe/PuuccshI2kP4R8RiIuXBXQtNvJpi3e1jOhOHD5kMPA431o+e6XC1ZbtUoLY5EQBfPtAWr
m7DuHD0pv7tvF8iaIS4D7f/CrRgbyIhdkRvsCXRexGKD2VC7Sdc8dWhqBCyHgqWb8Jl12hgvB6je
Vl4eZVUzVrGB4LJUstMV9G2f4Q35dk9F77qTdVck8WWyT9WaPTkwDN1RF7HjB3lEr+MotfAXqFZZ
129Fouw+7u5634Z4bBuZ6k4ct7EWGvjOMx/N1ZJih5hDLqTA02V8/0IoWkZGJB7V/eTP+/tgTAJt
HxicYlx6Xyrwbx+qqTmPl627vSXjcLQyHPvsMGhRg2UjBywgktyTR3CrM4ScUha87HrD4lJ025ZA
/ot/k1WS3v6+fcsnS1VtE6V63T0EGGE0KdEeuY0tyVx+cnrQKX9X5/MVEdZJaXyaoiIuu1mUYRRa
GXOouYOHDxJ8MCXZBGQD6TsMctlpF4zoYrUhFSs3bU9s9w0v0afL/O0u5WHXLqvlmVDSAI7gY503
bs9DlpWjZnfxl0Wqc/uJisaakIsrqwAj8ETbA9lWGUDF4sNa8+lpZq5jt/ABiKkhDYw0oDvLCJIg
NlfrFARzCs9ouBBQa5p9oBzNZrWOCEDob2mc4j3L2PZ3Ws7ys4IaPAQ7kB9f+v6Mf+aho84BQISo
rV6H2Ar+cA5FsgdtCG8CNpU3a5nVFg96mUgdc35//xywRrzZKnDEEiOC5Gui/CTaarffh5faXK/N
s4fn2v8nzzPhMVfe1nVbm4K9/VRFQv3EsLuq9WweaDymF+xzpgrpEaXYleus69jj7L5Di6NQBkBo
pD9BVhIOGnd0LruDQYjJUYq4KjZ8HSBjmRCgnus+BGhevOgJJTu/RY1xyVfCkQ5G4/a2w+Tt7JqT
sMnwfGAm8LFwQSax7q1IX3Uqg0jo7Xs/FING5eM0OllSiek1j8IVNsa+TOuvoMynQ2qGDcutqnu2
MUKrxaY/kTUmpFX5FLU3F6OLsWIUPnO+mSbPnhoC4DYgb7mD6aS8vKpDWqIF1tkr47GcAc8FeslP
iV1N7aivhJyOhhjcfnSqPg1w2h4YgKcsFs3VvcfmqtjAFv4//vD1O/VVUKD5Q+52CoDt8XrlL8FD
wgClapMN7+Yih9mDK+Vgj7BvCzlE2PwUHcda0W5x4+3iA0IYoyuQaioBODzS9M6R9bEuYQuQfxvx
BfBXshWG6l3FOTTW03rS/C1GU5472qeIT6goNoYn1uNBmt0U/S2rBKZTPb9YwPCiYUcMbrXE3EpT
VfkX168Y7US67aupi44pvpweLz55pwVrqARputXInVcHUzSzbqDHP+sPztzeUN8FNJbpVqF+VGNt
43crZ/f69JrJfWgtJSf+/uUjK5fib10Pd2uh1JzAaoEdrO02HytXqfEbysPbmzfO/m4YH6ovzbu9
8JToOxPIB9ElFCCgJQCPl4TAXJ3swiSKiXDgAt3JpdKjk3zeTFW4G36tia7jPoTaa+QYTWYSVY9h
jpaWoDECsfKiYnjBIFymOD2ajhHUpzaNpTfIVMkGc7GLnNCGlBHxxQcQoXN+WTho4iDrPYj24yk1
X+ldhtybNvnDrDMUJD1+KSW9EDtzj5LOUcUDalnwUOG4VhFe7/P2KeXXWDRBt6xX8h5kvlhX3QVf
irD1dAb+DpLnw2+ucMbrV6jyH+38dfTQQmPyhj/XWJwzoIYFkH2A/1oMxfmhA9J/8qJjH53DdP6S
XiVgsNuKIwj+wFuW3EyU0yByajyUh0lvtRTftXBdOLorlYUrQcHDbQMEi4W+rvZKJiHJivuTx0Qc
5+lXU4Qek+XiwB+UNKYq8vzccIYSwJ58Vcy3C4ywGBbEH4DQNklN9eXg7NogDO2eGUiCce7Aubz7
8RNmOSRW9iAbObfkVFYce/ISJo6fOx0u5Pt86VOlIpZrdmtyA4GEHUZSBSjMVQS+82gA+24rXHal
j0jHVwEu1wRPPTSOWuRvCodymxuT7v9c9ntr9Pi/hC2LCfSun2+D8gYhNCIPrVWQ0eRQ9wcF70Uv
JoZNn87jzb9YWZiRPxbx1rvO249XYl1fpj5entKbsUe2zKoxkAGB8e7teDJRsYp0hfpXUMOK66lG
TbEx4LRm2JGVG4HlEmziyW+PdD4a6cdDN8JZd3KBZyVp558NWMMSifsvtnMbvw3NS9aDzgApCUTD
FlxtAsZH41KwKKbjVGZVoNi1B2QBGB+ghea1UvzDfNFKVdS289Xzl2H4R4y5z9xVJ8w/SqqdncCQ
XDhURN9ljdjA1NI/0Uz2QPzXYyQf5eNFor9CdXJEnh/qlzMdXP+nZWYEjysDAX4r0HJruijIUAjB
TIgvdixw0qKlar8I+AmheVDOztZCblz9lviDUzV8JOkFegS9eTLqqv3x6KpACU83b8ifDypWeHY5
x2+mneKNFpKyF+C7vyVjYJFM4gFmy93yRttV/YYgLHH6svEIJ/Aikk2Z1yXRp+QSQTzRqCkXnFk8
kbf49uPj2aYk+FIACXFV1F9gvhh1fV6GCqWXCBRRk4vIpI1o7qjtpzL+/5TxMyjv0JZX3r4T4Bzx
Znxv3Wf0HgQLJm61LLnJqUM+2V9OlFRA6p4P6E+5jI2vtRwyu1jT/SWyyaBDB9eNIfq+s1/HWLY0
7LKln/+UMPZgcMgG9xi68kPTP5/KNGTJIKpSJxLjygk2oah4kbkPxWSEMdb7UhoaEF1goZchG30K
YsJi9V774e5eROhotrukt3wvPq0YkmH4on6sqxCNEfRS2Ly+mpsPyblhXm3PKjCxQUDojaSfwOxy
0QZw319gQwUADe/92Sh/cbI5Rikel/mG9t0ag3hfRf3PuIUHVnaOqbm+8+JKItFkTNDx1DOeg1u7
UyVpsQKK51eFrAc0IYVlxZMhPvv5JtwQdes16Dab9rMulcsT6ghhirW5F5fWAr1D8nOj2sUq6glk
HVy/V8Ww1h/YS+Xw2B292ZvYp5IWfzTxLXj3l7PPXUO62ZMux1SV1Cr0HLjND7Mn2f1CW5XwTF4a
fNZsU9/yD6RFD9HdEFPhklGnJGORxG8lKYOLhuZmxX2npTKtp406PNXTnopV/5Su3cttPdPMwfrn
3ziL4fZObo9Of6TUqE+5vuWICJnyWuufZlcKQ5mhSHNKtBS8/sEMUK3oCh6zT3kLQEwsCOg3EoB8
we8llZJ7h6B/JDYeZY+KiBG7S6BrkGvU511Fps5rOFIFzHlB0/KZvGVcpCmfyzMUduWR0uPG/TcI
hvx7mxfura539azKJGJQibmrMQkzkupsNYi0unihBPqQHU4YfljPsanFXs5/fF110slv4jdypuph
Crqs3StRwCud3DRi4O7ENM2I6uwNT4uFOcbgOc+Pb2+5rTdW75sGbyNPN/W99TvqNl+w7A6wugk9
L8ZKkqDYoOQO7yMmiLkDECiIyleQ0zVE/JXpbv51hpzoswYFuZJzt994ouEaMlwbSUyBfaZfdEr+
gXK4t8jDfUCA5OZAGDA5CwK2zjfip6xL1srWYcRI8bFDvTBnFwbWE8lUPVJaH8ZiHS6pgV0ezqQG
68a+OuGmZICPfVYiqA55KWP5amAfFNn5+9HtJjW24u+eUFxjefKKTyEjp2eYWBXByfOSnYXFcZTd
RHVN5tsfdEMCkSX/6hl/qiymZZMPWqtpG/YgqvfTfA8puS12TzwOBxM0LrbR+nTXrb+VQu1YQUNq
j5BwI4nxyVdjNomUjqg+hE7FgTXjunaD+4mcPDMH9epWPGnjEOGYltzZ94fzSumt+Ono5WbLw6m2
0TXXe8RjU5cQbZfB476Iripmw8cVprm8nbJFJZe9DVWTwxEgGpwMgMAsgGpF/h/Ew/Jgv7ic0v3K
GC2ZKgyV3cSs7EpH9nTfeyGuqTu4exHOPkvRPDBkJMwD1alVsbPpLe+xK7krTGswCBXQgLMqyinI
CBtoCBPVL0O7zpeJ3tBq6/y10azSXo1lDDYadO6VRgIjdnI0GW2Yi/Z+mk0DY9b4mednmvOdnNTi
BrzmcNcx1KhehHBlKa345lyDhfOI3jPiLeOenIf3848Sl72zZI6dcMmUSaWQCTEo3LaNeyOBnKt3
OVKKEHTpe/u8vj3OKpydN14MT6WcYFcz9z3BZK4CIYx4bnWT0zXZzrzsoGswTP9LhSTHoj7rjYUY
ahBbgXCkE9QKaZ8eSaqDCml64y8E69iXAE0rQGtHXWC7ZrWGnNrcx4qIk13G5ZZdjd0u7/s28HgC
kDAlwfCCZoD0JKbp5cu2Pkz0lN68QFezRnqrjQAdMngvNs6hhc4EsfllVyj/K5ODUoe1eiqi3tNY
lmpPdcgkxSD8brdKaPAVz1TjrPgIJiXEk0LZT6wniT7yYOqWw6/d7+GjuVNpId2MjGA0lV6eBhQy
XnSH0YY4Iv2+ivd9PpxQDtQbVO+yXPaV6OCLRTdgr2o+Us5584muAHBEv5blEE0KCksicEV2rKOE
5DFmRAd40XeDt+wJkgL4XCmi+i5izp72wfyogwfZlp6P5VM5HFzr8e0spetNgxNrBu2sADGbDtcc
yipNq2SsVYaCzH6ydVOg2UgprE9bA3SvobuuuzJgCMMooXV2eFqI3e+IUShkrR+bMFuRHF7sGAQR
axKTI0B8VujBetQAHipvwtwGJoES2FHouPcY2x+KnpmxqavSXy53OB2vaXncvzYRdFC5lbjQLI87
cpVWfPXH+5rISXnwqQ2bbH9kciGQOyioJJMZkrssClmEBLUlh/OrcEfxZONxHwdu8D6/mWqeBGrs
g0LoXGzc2D96Dtv6U2aZalsMcASEwjgCt92/jcMQglyCKBhDYThwdAKcxv6pSVV2/Ti5Urzz2hAi
o5VA961fzO1zfliYliZMdgVqPYjhqQtbEJw2mqfkI23fTWWqd+7kLR4618pJF701rSI6DPKp+cDB
nZt5gDH8sWTpJ/frpzUxAfsN7tPKEU9ac7se9Gmegc8pNr8AeRBv3wniFwcpoBHtBDqCbBWaCxtH
mQ88Okq+Xk+Wfarwq0i85r5SA67AhJCoOvXqXwXBFjcNjqAEk3PCVOwGK30wbD8rdryNIBM1ZVoJ
scWZ4WsQ3GGvMiOCY541hl6xy35Y2zb9TrTS7GbQ2ds9CR+xtghgrLYTlIO0CR0Jv0NoNBY/wQsa
zICSM1JZFMIgDY+EHHqI+BUy+GDTEHGHAwbHLJG9EBE6BL/9ygAmQb3SKsYvzKlOjNT0F02g0ggd
kPSIBuDLg0Z6VzM5+TbohE24twLvd/bd0kSvmpqSH6EpP6aVRAk1yeHUMcbZJ4TSBTaBPUfbLZzg
RlYO87ysiwDEz1yJkDm0bSKVaYrJqbN76bwVz6ad+Hg5dhJiL5Xz9kJUh5vhu/y5G9C38JfZ9oFd
TL+GGdpwX01QrcTRP/cQPmgMCjFfrGs3SOa+ZHYqGYuNu7iRzHTJmjWwC1x89YZKeumefqY1qXza
DB7GgwSq84z69GMzrFRdfBi/q2xCsCJaorVDJp3ttmgv3KqhCT9AItPiMeHokBcWvareRmLtriiB
6jzEEVBf5o6ghej5DRI4aRQR7X9cZ9QzfYpn4vZZl5RYAzkc49p0G0c1pwsFSmMN5mUxe0G7yfZS
iS9wsK43n/gGm/pRVePyu2otxiUtbguLmXSGbHPvtP7ZKFk/dSlJBSD2VOSS8WW/U5IYshE4rC0D
az7xFiG7vH566Bz4JZIllU6ZrYQE4ddzFk4dX5+X9AwcxsVt1L01r/j+wlny+/zvhZmY91P0CIYF
JfLaOfn9/TktXWCbEU/GPBaWodSQ9SSah/vXn61EtvN+rom41YMYUJeFvsTO0XaiPHWtKcoxcuS+
HALRLD9ksVINtANSSV5i7AhSjtSlbiQS9Q9gd3zjnazJmkkql9oXdtULcAkAe7Mo4JHCyFpfRfKh
46IPvnSnM6NPIqV3VPki6kcW+oH4+oVHFwj5+FnpNvYOcHXlgOCL+ScHM5ex1pW0kncc1GL7pxPE
eW4/Iv7k6eQZ42ocaHSFNelFoefg8zzR/VwXYaEukNQnf0TKJ3hYum7Yl6WIGx+6ZqAtIjv0ehsj
JW4PsB2HLZ+3QmlR2rPVEmdH/rO1y9lEX1/y5KkvwFmc1Es8a6GPSC96KoKWounFIX++yTzHSgsm
1xp5kKmHqqMczumr/aOiWa5lMD6z0GhZBMgM2kNpuz+yConRfo1cEfgZ8EboTVET4f7X0COYinA/
Ky3vkxt/3nXq6uNRcAjueSI5PizZpFQ0ecQQ25SgWWlvowrnfEDhE8A44wFiP6bF0c06qGzfzxHu
x5Dy+Y9MAm6Plj/Y0Q66uw2i0Iy8zgsPBc7VzVbYNEwPDjFGoKMEkrNZU2fD5mQE8vXB2MTvhnL6
QxL9HxmR9/YW6Vbmaev1JY04aF17GV4Rb6J49Bt6ryCSdrK9VQvzUByC+8/X7JqjypIeOf42li5Z
u1OWWrivrNVCVzZPVgOMOJmB+vZHqQlRdMn5Jrf88fky13ITmfHqBKulFH4N9HWzapbtby32DxhQ
chheW0Aqw6qJRAthC7ESqzANayEVerT+KerkmagnX08IpHQohFppuGrZmV3BVwrCvUQxV1/gbw3G
ScsA49pDa3+y+RZ25Sd4R5EjNFGmM7/OyaXs1Ck6XGCcSPRWi1tOHWIbhN0oiMIAxM84DfHKCv43
/fOnNiKaRg4hdaqR8FCEsCAF87qlH4NW9ZB/JdIriWMqmnXlNEw7AvG3b5MReL8jZziNgc8GkFp8
Sv1Uv5oQaaSCgwU/S1aHqIIlKNdji5iCN0IqvHY6EFhRMsC3EaabKHR1GWJg/T2ZvbofinNvGRWf
qkxhjyDik55mw02aJ8zz/U3VLmgipRU2hLJRfpYd0gYblVtIYw/h7kzwvYtGuLLqjUf4itdpChY1
5UPKF95UHH7wlOrS89RAqCmOBWOofpB+Nlv4Ek0zARvZr0YbyMAzFQRp+1GbKaiKmUibKRhLysUu
Jd43tCJWNMx5MQYzYg958l9Z9cv6NRcdyFGzSMU9TtKhLKQftLoe9pe4k9XHPJYzn8HT2EV4FyRe
iN4cmsM+EGKs0hpjfsxNMakU2ro4XVST+rcmQoFBb5lRFdh8fxyMsKvISfuoa1Xq8KHSmzKO3ovc
jw49uQUQnPSLz2Ff8Qc84nNSb+EBCxIxszHTNXhWT65Kflyt8fi7eU4aM85lytoHK0nXLujQz/en
/nTu5qDqZ2tU0tCAuZIQZT4Ohgd42ddEc2WbmeskjI772ZUySS/OrTAHdTgHJR0gMNerYs0vrMTD
RLNIYP8eBaxlI1OkkTXdwAYboWDgVAGCzLMCIa03uw/NCadXgv87Pq2BmGx8zixGwMmplzY0qmtT
dgb281F5ZqbaXtLZQ3yZSuKkKU8KtIL4XGJzTEyfcnDPw2UNeQgowy1dg+Ovt+KtUdjU5oQQzM5N
ctjs0zvLwS7o2UQ6Tb5zTApN6NmX/oeBsOFMv2okesxInb0pML0MpIC94khIy6qVggGqpp/YvF0V
/YuPVbMhAw+VpmVBr42EzWEiT7wRm2PoTind93EWvWsV96cwT3ik3xroRZ7zqnhtW0EglvLVGYxS
QNq+qZymg82FQxoS7VxsoiBZauELA2gjn1DLa8A/gZ75Gk3uu+/otTWJvl1HqqUhAqsZTY5I/kYC
0sT4lOgdQsv3c3St0yHzq8FWdFkxx4CjFMWAGpE2PD8GCJmd+tBmUJ+CjVeokAuC8VA3k6CuyyW/
H4oZH/dR8av3rfNwRl7IK6x0S/HjwWHdI+Jp3pfcYXrP8bqGBVyKwmwUWyHaiNG3VDut1UWxFLrH
gIx8OXGCOs1yoN/2/cKtKnCMeoBaZ4O7BNsJO0KxpySrbQIp+oFEBuCM5Vmo0KrXJ6snNpFl0s2L
zTJGGRXyaxG9gAvyFmlCJJos7SY2Y4anviDvKw0iIjn1uCiLfL/dFNQSDk6kjCbC8iD7eUVQykun
GJQHuLyVFLX4ps1zaXfHr2q03SmqfSxtgV5I2KXqaW/6Zx7yFqfF68i6dgA4pv5XdmTTm58Yszs0
UACqYDTHcVz76cz0QekGw+BWnhgcr5huSBh3TMz4V6FYmx4NZ5T2bbzYXJylykk81zBykg0hT/mH
/uTZLqTk3XWYkLm3BsKIMbUbfMP7SBMlHzUqKKjm2rewLfBuNqgjyc3JJCnzZHvYJaMRwO/fcJ8h
rTCwzkdEWROmwKW6clUfyfg+ilDZ2LzHn7iZ8bNsvy8+LcGsxGdirfszzGJ3Oul5+g/ke+yeZZ9g
jFWvXkS7C5ksi//bL31ptIJ4pU5kSi0z6ULYBI/Jh3ZbryxoF+G66nzGBGfZLk1TQ6swseCXAOaO
rOomJqimR7YywuZDB5irQ06qwRqYAsn2kVczpSm2L+UMv4+eJzrKEGxFQqG6KMefVb2KyXHYd8Wh
3fzwnrSe3UZnmt/VjckobLdoTe1PpbdJDdFOwiDgHavdvtwvWU7kayZvbFZxUhzsxYTDSpAIT3kS
ZF+F9H73QAHzQfz6o5MXZZ45rTV+7pOkD6QNQI44IlNwipSXwqHyIBwqW8ORI7yv//zvAkO6qGdO
veufZHNEKggw/0uYnsSBb/vpzSXT9NvlvGrR7nPpAq9YJuCnJpoHf+Y1zVfxmLyVqzfEsesaCD6c
9p/0FmXKfJLCzCob7ADgbHYvnr+t0F1Npwn8TIjBlVuUB05IyQvG7fHXj6zJyEauwKd8SMQfkRa/
eIx2Nfm7Nm/b1NkSELlVdiycZSU4eaeH/OcVLIYKhec/f2UUCSMuUOtx3TOKgnwEDMZ3R2rucbSr
j4WuOGUkejEOjw3CejJ0lOJsnPN+ywbegpGDn0OjOq0Ay9jBm0Hi4rwAQeqJXQYB4dZ6JoWI4rTW
KMF5IRRwCU3veUy+BgqqlhlufkoaEyZlvwu3ULl+lktUnibbWhDMS7JyIlSkTYmAQja+xwg/TDq6
oTAJj2umnx8676/JlTSgdqUIEQyU+Cf6v0ywbhPHed29itrytiVQaCKZdpktKfP/VZRi+61kIKul
xT4jiuU1OfR89ra5/5lti1ikTS5L4LE+k3T8lFvzqa1zqT+Cmp8cwD0zqZYyA0+RS6+xuTylg4Eq
ziVnat4tEnVPNL28LboWK9xSQPc61DRG1KED0gvKX9zZ9Px7KP7apZwmp+datLb1HP7t6PVCwptc
R8q2Eof2PtNVB7sia2UeKDreeYtQpw8MgHt/u40iLg1BWScIvETPG4yRz8490YVTBlGV8hCQQ1lw
eo5DCipnneYvv11NJKyGASFUfiLB0/QWWf4TYjHOYfojOvVtFkebG1CTbpWPdAsdmAuzJssVLj+w
6Gi2nD3rmdP/CJiOFOyE0VsH8kOXFtH+c4MpHtbTtRFX6t8vx8h9nfDXozXu7bVfw7Uf5vfR4iNC
7GjWwRpxV752sy+I+2aKJuPLzWCeWcnaHd6fX9/M/arQJFdPk2mx5JxIkbDQF/fC3kGlV8xCCL+4
HAgG8ZmxShmg1k++v2SZXQtzJ5UUOY3mrsRv1AZxQQRREJGe20X5AVrzXW8CE5UoEt9Ilt7pxEll
6JggFZDCrbaIAw5Uepsm1O5S3k7UKlR08cABngqoqj4+ZLF0IzdD3l680gvX7GNlVldTGgWZCjHh
XNYBGY5k3NiAivCwqx+f5TLb7Rl1D/QYZ/v0bTUVfcWoBWRk1Fpi1XM1hxtT0Gkc+J/AKUQz3iBQ
0PNaER4BNNZupAtf4CR5GVkq1gKFlPeSvYwYbNvsN82B1mbrug9tq8LShJ9683Ru7SKWTr5+fBBE
xTTikWcdxkzSfM/MvTqMxqkV6ip88y3qvIke5+yzMTam8ehUA0W7lXZxPYQThjoDxN8+X0HLeV0A
8pwori7kO6MVYeftOExgSJwIADDqlA3NInTREn3hVkQadgDpo/tIL3C0nyDYLWu5Er5qGSuxrHjj
Rgs2MMkUNnd4Xy502PBufSvJJsov5UUt38VNXF/fMitq5SWdO7XVOuHBq0mpuqzROmXpFzM/LxXk
1IcP5Y3QmqEeNfKjZ5NJdiKSVJWIrKSMQglufoUre/HueD5N0kS1/V15zJAB1viQhaScy6Ur/dr5
P3/DY5gGqKN2F6qpZu1PkKOi+hAc3IGZr0xMcGUZiRSeTF2TTTYEXhPopQSw2omXEOeDVx3+Fcqe
lsF2iZmy+QFA9edWZXdrbyYhXUUT/36+t6gzY6/lxTao405IpDFh+jHrzGdrwndxycbGwxQpGW2c
1hxtY8vpFBLZbOvoNa6RLbYHDU1FUgsS14daMk47PUBafVRpiBsTVYsZgfYc9Tl2lmftslbYgpgF
eom+QuchnsqT2nIaUUe/Fep9mQ0PQAIIwsiCYsyfj4xBL97rNemjDC7ZEv27WEGojDbkF4SXmrBu
Pw9CyBywJ8tbU26HToGgX8EuI6pO7uWzfCR+2ULKWBIkode1SKiYucQauuH5Uu9hjxpLyswND7wU
y02WfbyfH48lbfMtqh0CQRUY/N36/fU9ZNOrFKe/3ymBa7E2JHkscf+yADyPcvYQsxRy26WOLeQ+
v2rERGhdtJ4KhhXFM9n3FAWBfC5hhTER3bmfxx/Eea8uDgc/xTiU3OyXgpzekZmzeqhjREQpam82
Fn02iRvkCaigaOXMMbw/0mwJGzAc6Hp98mnczEKrq1aigIvEy3+VWeyxDWgvd+erM/61WlRLlmcD
VPe0OBW140iLLS+3r7RVGWlWGkGEWGfrgPDivvwJTqe5x6rV6s8njKCApUTLOStdvroGVdiIfDPQ
Z+JB81Xaue1uxvJ9NYCqJTJ+5as9F6T8nHJ2dpJ80k3bg0L6askCEmOHaL2rpN6tbvN6Xf8GDBcv
3+NZRkzYlPvFQ+c/DzQcBDPaxrJ3ke/8OpSxuhKBgNLZ+5Jq1WqzUOEvAZZDsD7NAlY0PsYAeDIH
EprDjx34jEVtRdV48ZCgoOfghr2bApFO3e6hteqWCIJ1QKqcUSrLn7PsEGfQeU5oBDT9YwkwiZh9
yU1Mw5sZAqy7/MEDoHZGMlFgToXVjPA99xbJaXgdLthHHJf812lT+EEXJ6LH6zGWJvnjlUy9Tl3h
HMvvSf5K68UbJivUwC0nMOQkTdm2TqtBOiyKTYQMwo9z6UYXgKBkLhHx/+vKzI5+4OXi5pfSUifW
ftpytPvMxbSy2MDkCvZlALzlXHdeDE1bpMlbFCkGyCzCb4ivuK44/Na01BVdOm0UkUAuh0BJ58WY
aozIXgzFsHXafAtXJxbl1XSBPt7kTPUdKAHRsu+3KYEfwNFZCMZbdYcyPdzXDEdEbTTvG5mLS7vh
RFusr6mXPUlvblc2ajBu0s/xjrxgA1XVuShX12aF9LvBP2r4mVrXkgyzFMl7C2kI/SGHhDXwV7P0
NlnhAmTFd6lwPAX5TiJCfvpDLijGwFygIcJi3/2rOSjm6nxj9kN2jkIr6cDY5ty26vnjksJ712WY
3gMj68IIpun3LB+YikhYAIQZdsqMEe6eUj7sEW0AMB6dSOfSdfLBVyao9O6DM2bb8WGa9zBkf161
Rx9GlEKaoanT/fcG8vsFL4Y9NeKpPUw96KdPToNttTi9F0+eRz/ql1H77F46pmPqPRn1YIt7IPy4
xHoEdLV86EamD923uJQ77LpsWoMdFDrVgzmFCbsjszclzD46XvU1R/yi8CoOAtxtpgqGtYyYjS5X
m5Jcjrs+lC8hdW3aruFNPUKI8YgUE4R5jyy8M3a/opvZAQCkBSUc5e7+MQL7YtRUVOBv2fT5kjqb
cSkygbjQlLA4ZD45Qm5ZP/+WRlTTyvsZCASsN5Bzey8pYfty9g5EZ4C0eUJMx38xwSBbSutX0bs2
wFdKfSVeSfEPCCN+MijpHPj45AQVqQfsgr1Zpw7+Sq/jaBD5Xz7bUaSW/JhaJ6dcrG6L2oYvOA64
sda8DzF9juGyOGmTzi+9Zg1SIy/ENAXLsOqakCBzo2sMrLanS/BwLFZybABNhcaeHUeF3peYekbl
d5TKkfspRqUgvf7qLma0mIN+JroLj2g+Dui8TvbU9tafHCilZIMe6G82MaNr5NaSk+ppjU7qzrtU
x26fSivgWeyUGT6nMY0SeOe6ITO8V9OoECd/V/AhQpUfFnsIRaNM/Y7gWq1W7OFX7un+6MznEq8e
lVYl2qJl6kxXydUbDwTUXAcc36DIIDxxrZ0OQKOjDGXZjtA4sxK1qBzzgeHp00akGrsc/9/RYmKb
/uRgHzbIur25lSK8Ma3aUNEnmHRhhQgqB9qRVHk0pnDoeolUhBVFcPW9B7WPitjDWV0Z0M9bqS+y
9Frt9yvG09ln/OBFJvpjZegnFhNGTBAWKxLPr91MtIm0Y8PcTsH1jrnxz35n1C9AJ85KWw1hqDlp
VBAXIRjNOzURAgB7xqPBgojH2c3g//8RQmoIgYuLZMfFPpJx0h2kGiG1ovb2rlEtLh/DUzIgrHKW
5FloOU3daN9GbVUErG8YrjVztsZN8sKXZn0CnqiJnFw+Ei4iWaS4wL91ZhMlhsEjtV5vO37urZIl
vR5oaNAweslXhtf5LSDwxR+WWPo2F6H0Lv9rVeoMbhlTRqrQrE5w1dSxHb8MnbF7/IAX4ARZ7h1g
4kUVgR96AVn9ziKKRJTMPpK+deAYbakhg7IsemiwwMVCoOIf8qgTKvRhmVH+y+WvfI3J44FJxCsZ
wJ/RQHQU0e8EIBUduAGmQhOymnwc6LDkHo7m6JJs2HA2i1f2BZSaa+vP/d1rMqHgUE+ih4ojgR32
DbrBqEeufbXFx/tDsDkKZo7waPvlxzeXGTyVMfn47NTMHhnFbUxQnwfIsg6y0RBcOUJipg5QiFNW
7GHga8tjtLYr8HZUmtmL9scGJxyFMX4OQeCQkwT0FzUHVijoX3BZeckAsFSf3XEmzX+SvgMYLA2l
TPBGhZZaC3FmEXfm+Da0+2rySH/lPhm18ZDHqpmmeyfW1fGCGf45PawBjrxf0B3Qb8iMRnnBaiuw
dWy8AeW2Gfo9O3hL9k/sSiH95bgm/sjXDXViuIjaa3zcizSRQuRWAzvYbgwjbmLK+zDl0NJVr8ST
KpbklrFWPjSu1xo9+A22XJosWY19jGDD/OqwVUtKQXga6liW9PQRZE2DLFTgAvhcAlDMjS1MlXWp
maeo7sCBedcE/TLyYt7fZVKk2K+jtkx5Fwu9X5rqnmt2dn4n4mSCa3KVeJlmTwpPmdtU+57tAa23
llMtWpyubTTzl7TVWqzp26w8VVNEwnS2TdHm+ZiJVLYcjNafdZW4s1TJN6HFEUSs3as79vLMjmpr
dq/R3KVEP+3LCdc9l8yYDQHtA0ZNeoj681VvnsF6Hz0vesTOSQ70efyeLulxEGRcoU+vtWbCJcCl
v3We/YaqmJVWibk82wTdY/7mtEfNh3NRrSlDZnu1pGxUtsmdtTh89IMkOPzsLuJnyCHYZMhv0mHq
tM2SsQlN17ZJUq8ktyr5F54XAUr4wdwtpYt31neqKkMYx6kQBjYlNBhGkdlFXFGN28a02v7gLPBx
qHXiDoUdGwaTh7uZMFaBf/qcOvMDMMydrdCjat81DlDj8jLwUHMT+c85S6cJDL1NkDYRnAWbJHJr
6a95JdkB/mw7DTjqDIUyQ6J50MKiqA1PMB0jJwnWNF2ZfQJuUTITwPFtZSYk7hi4C6RUrkXkrYGh
/lx798QUvwPIUZIuJqReCzUU+It7W8zwWPkbpuZv3w6DtmkEwgkCfMCfhHzdnpkJe9zbyJK1tMfL
6fxuYq4Et2Bi5OaI7/LLqkAUUyZ5paQUq5v/5ltXRqliQRsD7szSsa3QmR90Z2NtNRlShSdCPcvd
SgoBPRJ83kFxOYpS/009WzhIVQGyUHrThv2g8Ixz/zhMrAbemlZZdU9Fi5OHB2bwUasyndxqMcbC
JjtQxtkcRbA/Zd0zT9quxMnVZTlVExSfvukG3qEg03TDCXIbHmKlUa+PU37o1+DHyqddnhDe/6Jj
Y/H87THFyBNQHjaIntrqp1s404B7YOB2yyvvgX2zBY/eB30dKNcYZNVKfczu1EyDBnuNuhX8UAmQ
CRoCkgqYyexiBqQloRUleLrhCmQK2JlbTHFYjGMPDEOLrYYjWa7sJmPcQQ5LORQSCYjQlkV7sjKs
wOZnOa7jsf0nd4A8NFqqbjixfgPFUlelVVB+ugxkOSJO1m2AmIoJuWABcWFDlbhhf+qaGER/l28C
dBN8EvR8fWLb7mJJB2Yi+C/30Vt7zfUvUvIsjsHTdRzx3cLPuoq5oPDaRDUQ9TgrVDaaDUJ05iqt
lJq/7UdYhIiAewbAZEu/DEiCwAEsIVMvu6T7aJt5C53uayrTg7dQbiOhNIZAchsNEfOiwFSTGox1
WuZ+EekFe5BAQ1XMEIH+2s4apMsu5xmFKfF/aDZGsP+cwTy3qIughwyvXIxpESzn1rMm4GBxnVgR
a9Xdrs5GMtUb/qR/SxxIvDKCk4Cbwbxx64cRLbulCaVsUxQXJ5CN1mT7Mb+6YVAF33BtkkDC8bs4
65nv6WiqiKn7wHQMDfAmMDOyN4ZVn5lXgSf639awzl/rseJEOaL9f45x3eVXEZSnqV4ozQVAfaKk
C8gRTbQcJ08B9iUbrmrlBBLARDnoxcA1l89viinibskwNA++/GJoL4O2wTShrIV4lYnl+C6LkuF7
8nKfUGmlKWKxwnR4Lv62oljaHmTBP13vSnqsP6M3HuwU+GduYxl3ljqfSGkxEx9Yfo7kE0XjXmc1
y0Jc+lKVyAPLw5gSzd6pprtZzGpoxkICcCxFWn3QOzf7QeLwmNwoPnw+58Uo3bSlD56PekPh0M8F
2ZDc9ah72QrRyrQZWGXZ3LFFWSn8cYdcPikvf0mrX+9tvRuRMT3McsYFy+EzmET6o4iATgz9ggXa
sMne4g8O89JQsa4DYBmn0Q5HiSFXqogFhtNROfbALeT4ZyBTDkXKH13YevnVVHWHaFXwIS428xb4
dromWTVqZsj6rtCmsdFkHEonXFTtaEckH7fCOvePmcivfecjHpfBayQTxtCXby7khW2BN7VYNeDH
USnFTkO8nytvFeG98fYpeWdxVPYW5h2CZNr4SLPGVv6j5lXWy/G3yQgAct8xegsq8cESyKq9iUWJ
pl6lbQvGTr39jeSshq6vC1cb/CcK5Ru1PL4iV3WCl7hCjSFpeHos6fQFNRZ4IP0jHpVZORyVB2px
0nMrLVWLXH3AXcjYrmat7sagHKVSv7Rs5IbPf7OxUF4SEa7vQP/s9YBMhPH2NV6I4nV+xicrVazf
CQwboVye/Ny7Vn0bT1PYoEyZiWzXatuq665JJwaCcer6Rwl3azdQ1IKENKzpBhZOuDm90Y9mTG6t
wNriVhv26baI6EVTYDN/pBNDJWkmKXIMntXbBKNad8IZiZ8IKfzr9f4oOZwvKyXKsCDBIHwlJqUR
9+Cre3jDQq+6fO6qlVMUMM3eog+U/WQF+R2S+cYQIdj2TbbSq+ZK+osKppM+HWWZNzpvKVE6DDM8
u3k51ILuMK7rzJwS6RK/qmJPnIISoqpaHDs0MI5F/iyO3oZyu/uB3MEsyWlWSqmfBtSxXmndUCZR
9MXZ0TU9vr+798VGQlBQtyeusSKzW5eSZvcfX/UBLWTtmuDXPU6U/hPgV/pDKn+UMY1QPiRUsXf1
es06+51/llIQUwl0E81H9KOFZQILq1O7+wFUc6799hH1zGWJddH2sU2tH/tuqUgkPInXQJF/OyA4
+koroZ7eY355szKwKKJjLGKFGlY5LFAG9uSddiE6KHyTsURqmE9xWwECpLgjYF7bppP0N4PFSPwD
Z37+1PrhkzR20DryLHJyc7dudxzDIPJk/D8FnV7K7wbP6vkgCydkFnCJlQW9Mkafy47djYz/rIAk
DBoA5o3zRtQjGwRZ1oe8p5ZGk2tK/AUqpV8FZ9ukA3GH1IEvyoX0HiWM5uqEOSJePOod3CbXKRmm
H+eNf22pE99yWTSpbW3rv3UFS6UZE0fmMlkFFifouybQy9ZpT0lodqNDB1KKHArWy1LavimNN6kw
Bd/a6k3GAi5QBFmsvHvnNZsmFHpZYJcghV4zUR7LlLT2h2BpAvYLcGNYEpGq1mthpUtpsysQCvYp
+CmvnWNkgQ8BqzRnvm+Klj2bpm/+q9sfrGPsMf+plT5gMwaxQYi3eHqsAI697jL8SYbQC+RbA5oa
oOs3gRYbFcDSgblW6ArRblFXgp7Z1PY6OXegbEgcPRpmqWYRAogKEppbjQSLmeVD7Vjq8U3GnJN2
9AgVpEvXDbSAZ8v4w9ErgZlyr/hFsZTBaN/SEyZyUrq56HKUjyRFiesi+mdMO9JJdNpp0cf5T2TA
rWJusmQhwGIYa8pY8awGx0UJpFoZ7MPJbDynt9Lk4Lf1MuUa1eoy1b8V8pDmgObTOzrae5lf2sfR
fWDJTS85waYlzCinTKOMLRcftopCguywnmtHQypICJ4arWknLSacU1KcW904A7MMpTq6eNJKxehx
avf3+JhSmXv1puM9dMKrSUDebk5pUwTc75MNXapalThL5U6FlgNVwBEPCdEeyFkjQZPFJfy/wm/r
ZCkKk2KLPG8jij+7EO3aAdWJYy9FDxkPksW2F+nnUSJwcKT7WjQ2s092+pGGHp6sq28x7sVIcyfI
hSWsWZsRZwZsLaLcrEcwwuIubERwDlPvUbffcgvRvLL733v4a2D0yYxY2hAJizWv4JQpoj6mvlUZ
fm1F3+XDci/Bm+3jQ2ops6jExd6hfZaiCfckJN7LvIZVODEin6FMc82qhzPhg4fHnkyGUhspCb08
bbwX/ysSIUdBNV5amuMrDAQpaN5rwf23NFD4qmlV++OZPNUnLPzvoWX1SagQe3lNp8rpLOLpdOAy
SCQeGG5/zYG/6Y0+ju8BPDoPbjYu0/AN53RGg1D9IB1ARidqVBx/+qdNAmxjF9KggLY0qtNTLeM3
l/vVaGlD/a73p31yjFccpM9s0NS7ki/5SDb5KmYcgqemJ9kBeUfXcU9ZS1P/EyuXnZowrwIti/AA
MCq+W4Y8WngL1bysm5PUvj78z+1y5smiTqBZ7SgyYBGXrLXMBchyZ7LSY69+HqnITGc3RvENjjd0
MdZ6G4KKf6BZLJsz6CA+MeW2y5WYV5E0ERmNac7w8OCz4pO+tUmHH7BccJpPhCCkW1bKq7eT45yq
JZnevu6XgqqEIW91Y/IELHdtxmDyRoV4pPUqg4ls9sPLDc6qwR2MXQnQP1dnTjMSKOq1wst3SZXy
xRQlPzaBAH53cRuxojRK0+7pOoSNWJiwujRb8RZrOGdAw2jAHRFJJVEexd9692FV79bzaEEiviTG
1ttEaGTyU3NpMrvW6P/cx6EcdGUME2bBRn81OAdOlGikrEFXY3iFM8sWKRaGumeW01yw03UvPiQn
TSNHxfpDN+xeZPRs2Qa/Z1L3Wu2WYujnvqPKKmwC5lWeCXA6YClzqWQsgPg0lntfIbcZWEHj4UqA
sW8jVFOGXLZrXSmsy/8VfCiaerLPjNJBNnSFjAIpMVlJScxNlGTv0a64LB9cC1UqSg/cu4NalK0D
Yn8qEPbBboRtJQ5tqKzTsLn+2vn9rk9mFnKRr5uYJ6DLBY2T9/7nGocErjDSrgOKbcyx1prH5peQ
79czGQjIQxYXohpgEqY4p0ymJ7H2pGslwxLuUV+FlPV/Aq91KaPSQjPCMrJhbezmi4dHrRlTyZp8
YK2Uxc7IOXVrrQWRCcHqQmhszVFIRhYQcmmXTEDSYdlzyT52pUlXBAlqWLHl54dxGsFGqgn9sGCV
0LeVK80yJm/dU18MYwTMu7b9W6NvqutXSNCqDlXeOI/gJDxwiq5UnJ9IzRho04EEl7iv8fGi/tFl
0sJoLE9nfSAbn9ankvC12iGOMyeUjDpeRR1u7fmqISaYrGj5LzkxRednZgqFuMfVp7geKuP1Anyb
GIJBruYi7N9ErUtDM2pDv/KZ4TGAMkzP68LzjZg9oltd/eozJjKAgl1O5IVFIv4/cSSPiLmmPwcr
hSnoARenhRVVK1r6AQMtjmdDn0cB7p3ENNJHtdWwQ5JspFc+i4ZIUoNtykrk61R70LKUcre7X+cn
zO4ZIk41cA1w3CglJ0z73QP3ZrsXdcFVlvlmCVS299koz0EftmEcu65VlPp5J4LP3bIX55+m3xUL
7v/f7pVSVaBjUKxlYpKT7BdSjKdr95v8vgqDD19fYpCXkJ5uREq8N5tBeTtpnMoUQu0r1pzsd9au
dYKuWlcZA8FOZJ1dPG7a7wG4n7p9kOHktUdP9TzBgJsRc7q5CAk91M0twUgM+zDMBvqH/7IE2J9a
D7th6NS2cIJ49bonY3PtrpYiClgJhrjZZx8LXuJbR1jSfQkyXu+TW6njulNYVCYgORDsYceWk73o
rY35K669sQ7UsGFGO147gAM8y5OYiEb3qcQrmzD4UKigYcTtp4swtDRxCoJSlwDmmlkau1d8lAqG
oyi/gyn2XUjKpMkDjHBeZ71T2fo5ojHgKOrsd1TqvPj34KLHG9/Fa0cy8Bul5ZXUoQMFUUToGrgg
aVWYljQ0zWQrpCUnB3RVfy5fzVJfdwTOW0GOfepBZ0hKyK9UGkNV7NAM9KUecOFltlQc21OJ/zju
9nBDR6S3Gcj4gAcq6EeQAKIRSj4rNcuvsoUprV1NiEvKQ7ZCwjgHO2p6ldMHn8stQoRLGmPKMTqG
WLvN85HPAn+hs66zpdfhoNsLY4G8UxhajF5kB7D8PIHTsn9Nd1NzEcKVNfmVQeHxwuumf3+z8TU6
+2AgmFAUf4RH8NrZbAfwPAYp+CBn7Hw6rnW/I8T367urxplpvYLMqYqjVVutqo7V70oImgsPfWgY
OF4FIPfFh2PZveYhkC4xb57asCG9J7zPS85ShrYhJGSi+oMzrBzhpokDk+4NIjwEZ7QBj/8aP2rx
OilmGBnE32Vkr1Z135PuQfgl7gGxjKXA9+rw+E55dv7zpe8Oew/s9n3Tw8y5E+ef6DWC6vmVYJf+
Ud/sv/sB7GzTrZ2pywqEQBc6FLkP5nfqAhh4XGsEuMz0Shdr6o3WZoZp5ZH7K5z18yiE0+dm3uAY
UiA5BClQGa/ib9LXp1S0G1oMKYnJnsHkM/PkmwSKL/f4ou5fXRg6XHozLxsFILJhm7TY6+pw4Xz1
XFX+HNMvJ1lwmhWQfMrl/5OiWMQReRN7eREzOcR0kGFFQmrtRNP7zNqiTf2tOqqxK03V/Qajx8Zz
PGz+ZpfTA1UcLZCRaNgI2lp9oF3W5Zk8EqU14F2SPX6FqzV3fDEZRmuXAMIUVTkdivf2hzsg0UpL
us/X2UkXfdgnFZse/QfD4HL6gA7PF7ZDVbc1YJDTYQ0hPAJEPLjph3wwl4XvWHmleL1SCEvhpHDS
no1cvXTTuzepw2sQxqhOEqi9w3AIo0U8w2nVdGeOAh5q5Qqg/0jj957pZB67Kt7cnf5D0yciowMC
ATGdp4sH7+0WtI4Pr++MJQ49GCfS2JzazbhpwUbzUuhfI4uKXPit7cr9rgjcbcsv1TR62Xv67cgY
u4e9SWTdYzjTRf+IDjwAoIEroe5BmVlZWZK56/fSjruxSiwFuVsZCFcBYbj0kLh0RMYm6Hxb+jgS
9BFheYV0qAEmLtX0T83mdSiwV+hGrvwhWcpZjAZBH3uk0J1fSUIMl0znyhCFejBglvsx7eeN8YpS
wPEV/R7Zj+1lDOrRG8Hl9FY2LqvrrCKwHdiS+0KR2Wv8ZRAYQKfVR0mdWo8GrC8faoYjtVG+7y4P
JtKg4P0zsglSG28sH+yD78botJq1f7JlIfFBtPdehT6rE13w0BhGLXYOsXGyZxhsqHa1RI6p3/Gm
aVJ0jD+C+xFZSNDbfB1ByOdiL6nnkOoTAgUPL7Ra9cmDLsuw9V+3FJjlrUFBeRK/pcm+bb9hxdIk
WcIMwbJ2ApJnVzKKH/9cVHfOem7kPPVjgk8nrNsdgfELySmoPYhLhgfKmYO4Q0nFNEV23AchCCTw
qgcsXh9ASHKwkeTzim6J4T6phXJmR2THLVNxn/U1mBEm1tXYqbCN2dxMpdCnpXrPwxPT6QSPneHL
xRVblY6eGU9QhPMgw/YeISFqWmw/RXJQxEl7JzOh6Op0Xhf5cOOaOwrCXZ9Fca5qKV/8gwQ96jDI
12QXhf32dLRO7TiTsKxBBN+UcYjvD/FFgQmUBqicJZFFmUO7uY0A4sd0uO0zksCCsScnvlbZ1qOl
Zb7vajDQrCkMrjlg+n57yMRHU7l/r6riFMBugPeCeyOMEqyOWLGZFSSoA0qfjYEKZi6wgU0hyUtt
+fMih/heqEl4QfVo/fWdBtPO+wjR0PbKOI/rPQY1mAIVuGuVdg7fXJ5o9U1FBCj9CCe8a7cMXvo9
JJi6vqHygr6CaC2BrRSHH86IxP3qqThmqXgf23JkkDA/CvGVU21EuklAfCSQOpqWmG7yg2abRGSq
M6yPjYnlSVWZASUwWFq5fyNE5Em7BOAxgY+kMRDDOJJmKdJ36yLehyrhRifLGnLhpVabxOUtmwvM
XtIZSkh27TNyNmJdk0pk7P0OvzC1nXmosW3/m8eFj9lY5A/RGZW+aAK8sKCKNqF4YDigGkOLQFUl
5Kc69Ry7s94lIRXnTZSwXDQihmdeBwDs5LOARMp8L2y4BITYqHQBG9FAZv+I4vgQ2jznukwcDjnO
kApS/0EJA2U1tlgOaemLXwZjmx08Y/JYjlqzPCJxfI+DDW0Li0WczzID2Y/Y4GlChdoV3+/pBslC
98nBu2/zYFdXz1K/1mImb4kk0+qnJRb4IVk7pvhB2Bh5gq3EE4fJ/gPM4lavWWVrGQAYcFutypms
87DPEP1aV2W1XSg0nqhjR0TxvvQKy8JfRYAHlWif2k1ONlYOKykHU/4L8DzTEMmOYg1bo0PuaxCB
o6rYInZqEHxGOaNo/aO4pAqDochxrIDqmnxS8j0uiLH0ly1OKxYemGed0DkdOB0AcIpAEfgUjGss
mGWP/3umI1eh4OFLEMgWMKyUTDeMy6HuerJ8OL9ra2EUt8bJZn+CXFEW9hlLpl4JzW6F8p6zspCt
J45lX9r/xu6itr6fh3afifEMVgvUGSVrjjNjShuOjOOoAdqeQD89VX5GfFRi2l5TY+z3RZFW1k2G
o21z1RVN82ydfmx8pPRq60vDCQIWCmcH4r2jS62yPs3ZSLggI3WiL3e9GZn7fNWBTboOc0zl0AJ7
4dSkR9V5cHh6qFcBbfh9XO6aLWom+zYMgf5mrtAC0xOCQbO0xd5okbbLSUk7B9cWDIhtL6FFGHxk
7A776jHkxwfkGwBUGv3fgCWx+02A9rPgwZYDH7xEfpQJ6pX2bQLANEEP3bjbsH0FmrKismDqtEqh
t5qj3NsKAjQobtfjcVxskGm4OJjuoLz9PHVG98kheHIosX9scgGQ8ojewrJQRistV1pdNuEfXXB+
mPFMsOK3xV798SXdR50sx6FJ4jClt92GyjPTBEbROagG5KEiL2Wnck5Eq+hIGifzj02cJqxP8npo
KzIyXnqrdzZosXkWcD67/sEU/imh5igPff6daLtA9WXuJU/vIFMR+SVCBpK9+kDngAkqNxrJvpAG
IiFayCQZ912ZZJCq06pzcxe6LWENrGo22f7LS6N/tg0QtSFAZ+598lbiV6aY8nOnMP2qW3Ni4agE
CMJqRFwtLuhLbn3kuVYMya14wP2N2MXpjWJgkfWgxwKHqqUPfNFmydUATyusix2MQknfcnc74gcr
zmd+25bGv1oijAxIoR1OLDSp0CLv8NrXribpxvy5JdtIpcGmuDla/eDlbk32HHDEHGSLT1kH15ph
BFWGTtPOVzxwY3Lea8Dk4678uMouAT2GkI72tRGlrtDLoYQkBLlJ8WI01BCaL4OUdtxl5YmzuGfB
pwkWMbsxYuNiepVM0I66GbE2XSr/mBGpLfjLgGjB6wElSe7S6LoCuuCjjisHbDbouw34fYShCH+i
S92qxZ91jsaeOCWKU2DDLBCY5u87JYH+IZITNuArg4QmttKqHQT9we62O70Kg0u9PLefvPhrsN2Z
Xo+ihUrB2kzgIp3JsjFlNb4OlS/LX0cjarRMOCHZ0LfY1fFMDk9SE8eO2VYOTGlPO1fjAaC3wXl9
exw1hMNukfbLSXlmTsphcqFG1y5vQdXRhXANWqfnEyEn8MglzpuDKyjem5aDm1/JEc3hJG1yVbK9
p2e+ckJZqy86kO61cbIcq2zCmXZ6oX2UG25g+9EVfpkA68DRTXlXliz2HHzh56G2BJY0AaCOSQIY
WyICvy+4ROBwadrnuYshwtAV14etf3vU4M3UJao2YLiU9KL/64aH+twEWFhFZvID2gxXSPGrxMB3
b9s+Ib5LLrpmKcUMYbuH321kqIpBEicWGHUprCeChC5P8DoJkdyANryaG3N7T+nV9qMRfENL5+Vv
AgDLOfKu9iqT9hOs7npkLnjxioR/VZhH7B3u9KUvr9KDZy4EfIUKHL03frZH95G+ZC9xZ1l/S7pB
4psi7z998W9JBteiixDN5TuajbMfuEdXfkjxs9oDtY4BtLs3JXIeaXUsV6gq2G6b8v1neTHUBpZH
kYUMozaHevjXea5d5IBBJXLv8IwJ4k1sAIF/md1nRClbTGWwQgXpGQQr3WYODLFYUNUzEGjtvfTS
7I1naHmEJMr81YRe/FrZtuLcGqYj3dHueS0ikImMaK9S5gVfQ/YmHTBzDzJ+W2g1XbcWUFdRtbqc
y+KmLorjF0Df2BcztOgeh8DVnOVYpUcFqGn3bzgG5641IMNzT+flf8wnhK8KSRi91ODZYStRfS4A
xF0ELUuciUuzkiT0rZ0OtA9SPcEe0hfahGNOZCUAqdeJ0JA9L5QsF72ZlDjEHZUMijk3CXDI23qS
1lnrKSZu8Rh8nGIjec+cW0F2gOlq8TSQuvMEvOz/lcyGyMOR8BGh66jdNGOHupPbvKqTf1+3Ht2i
rzIAD/onh0C3MTFBPDwQ9suv+eID6MvACHH9EII6mH9qpoVn6SLXP50+cxclHveS+8qfW3f/i3BC
TWnc6A5ZjRL57nFmybEMHYAWJNr13NEscmcW520/W3TlaYLYOLgDWu0My9Ou0x4WWG6SdtR4BWj0
FJ3Iw0is9672oSjmYdUKhXsQD0wxkXKQedOE2eCzO94vSZG6sgT++mLwxGntGfxMOdRlq5z7M7J9
N6jisSQxPkFzrr0WuCm6s9ocj8WN5znqla9Q1uH8igWVNFhP0QC/7ROMGIG8rcaYEVKrxMfIXCXP
9gjBkmkE73sp12fVIKVUYXTBYKVqix//RxhifUj8pQ1IrHC1qMJMh0xNXx1TkDL0UzkEPGnxjecm
Vh9rMBX0OEHWQ5x2yjqfCvazmz0PJZ7QXxoFx3NDkbhRaLeS2l+9m7+MC70lYoeDqChfq1qYPI8G
ZnWV8qQNEuOYgMzF6ddsrSpUAtQrbSqJI6W2m4C3YPl6+eCEGjk5R61UYdLeAIKZ/VtRTrZOagqr
BXrApp1FatXjOQXt+akzyf+TjWz1loqf1LuTJXUkJTveUMN/H0u7/NyAg23nGzl5Dc/kADGf2gjm
9fgaphB1sEHT/LW8TeGFAsoZS8dcXKXYD6XrHUB2E7a2ZaBUYoA8hMna+a55yOlrFP7Uf3v6maJ6
qkcjq8GLa5zduMoDo5hV586ZSBPgBLksCuscpIguPqYmUInj0KWQocGbKWeJhMCilODnEsyH+Aj6
JvWmrH64LAd8oJtIMpYPu/Nx93Oq3cMHu43sIbGJDPobT/jdY2p6Tg99eE9If5s/1k4fImahvK0v
D+NFoSiyklsGHLypxzIKVnc8QkUva99q1Q8/DQjJ/j7DeO7imXXqqOOGm2vB+0iapO+ZlIv4LBiF
qPk8oiSQRUj2X0dOHtAeAjUfJ87u2g71UYVgQiggQTYjG5Nux+LDB+4Qlpy0NcBOxz/94Q46356w
T+n2Ldixe+H/tWvZF1IfzPE7wAF6GqH+/IQE2ea9/3e0XDH58peBAAahqTpCg4XkG97+TDaB+0Ee
75Bn4BbmNJkx0awOTQCE6GqrWTOUmNaHxnaIAITOrbdQLrdMxC+ourA6hB50M4C7Rr7/y9Enxox3
ghY8HePnNAwWSGAh02z0Nz2LLUw1izfyURsE2NnH1ZmSoJu5psprbC7Vx/Yv8dtgEHFJbxzmm1qG
V+yJhEAr0KDa0JLt5tY0GSxM0MKntrnBFB/hID+d6s9pVbY47zXQdFJ09xskBPizhis8jM/nIrDt
6bKFLbAvZ5I0l8JZ75eJhGYhU9HdMR/zsojp/PQxRPaH7jmWwmDj+tTzSluAXtFQIIocDJj4tusT
H8vjwCojFhzq07/45jUTrP+nNSnlu48hpnDLZQXiE25d+5HEs7NWBxFo5sNTjcfNZxlIomkOoowj
z3VnhzyqBjdfAdab7VQ3PcoaAC51Kd8J2ecAbEbdtsBtmXtSrgeXAR0tqz2zTXBIUWdgjngKuvYD
898LoxuJPPzx+ilNhEwySJoQGrn+opnru2Sv5iMiACYtmKeqUZLUn+hjYVeOQeRzX/cpIK8+GfHR
iZYVOxO3fZ1JXsOpX865Bar4Y5fVD93O0vlia6jlU5Iiaruku/XLo2/ud7QU2Xcwejs3NSpSw0aB
VYyH09MkPs2Ks4XYcbbPVceyU0ymU0WjHVmBaXIVkGfe5UTEcD/CMAYZUxpWHPEZPxNz7UslWDL6
JTsvYhBj51oOiB/rNr7X7fBC7dE525jjaFSmB85GtAkk954Ahv/eJrpgY3Sc72fpTLjbTzBaKpxV
3LMPQaHy3T4FSmUaiRVtZPIz7yermZCabTse5FMpiksnY8Q0aQN0/IA5qYzUp9DGVcEtFehgvqQ2
8l1MCHK/cd3CxUEpAgr0feBvus9xmY4vDA5JAxbFkBFQDpZxWuiSCvjekFspsSrBB6eZj/FZkRmR
q3Dri+oRru5hgd80uz5RYL5E9PpYQTHvZlSLMUxY6fDoFJFeDJpjZB/Kt8A7nDS2q4me1yjslPRC
msziV09zDAZFFoBVsaeRpGCtVqWxL+Mjgh4henXgDKaL0Q4gUDOwSALt9/vTGwOWuxQ4SNT3yfWN
rlcpnmybuGMy0cWk9bkPqCyfQGZMqwIcudgKr1SVx/Ht+DR00BBEtp6Kc2y6Yts7ijla7FMj+y4Y
UUvXfTXsWSCxK2txiabtTLKTmBt3T0IE+mJl0BpNhCZogTfcQG9QM/m8bb+HuoaYHHzigNUqXh8V
fS5qoW/xMLNn1Ms3xWmdY8bff3LWPTRKWte2dtpM37Mz2aLRW9prNq94Sj7VsWZcIl48mgXxZ1au
6e/LOJGFZ7Grt8flC3kSNim48c0KcEphDjBWPu3w8hgWI89fkWDm36Qo7ckLvrdIIcUF0UDqv+tg
uIY41upXtiWFmcb+4TL4BU1cOsxj1mXes5pjKFLfY6iP5vS5PXyMmvbnhTf5zrlaHtOS3/9hB7o1
tMrMupj/DY7tMTUCoNhKqLmQ8/r9OtvJZ7LnjpJhHFPml0hDUtx9F1jtrmqsj0Lnr9GbowRu8XzZ
Ix9qBhvEYgMZVo9HHzBhkHf6NFJY+oqctp+Xpwrq9PW17PYGpv0jwmMlV+jzyDFmSql172KbMAMU
BVOrZ0FaYFwPHSnbxTMHC6m1sGDAz0+um5UR3d2co50ln/a0bvd/0MtwmxNHuwMBOG2eZuRdcwqN
MHDvrqPjNgjkoHb1lYBTNRRt+6QCBUlNjiD6luY/L/OW9CBemOG8cET0JJ/I2iwAyk++dGK/v0t1
fkQPnb30X9rYqfvv4QbBYWmotoNrnu2/bF7VDuDGr/moQ9jZXr69Bbqobki7N24gBBp5QsFKIEaZ
QlnkVFB7KCBF3DIGFm8CyyxGGS6g7yTq/UiS9n96lF948uroXAcpHEFewp13tJoeU5skhFAi4vol
w/v65VnkChK/8tFgAIQ40iwBjbhsyB/24aHbqPmpRNmPTJZgfLTzrOToYMd/j0nhw67LZ68DDZpH
urUnV53pe593aGceNjns6huxdqxeTXGs8C+guNqb+WFTCgdj/x9lA1oC6jSowHaxm3dNvUMdvD6k
HPsmGqBZaW71XJPzd2/Jy2kgGTjTbLKnE+eFs8WQpUOBDMslmHBbFQSLh9fchSagd1d2rwUV7huN
SirdGWoKf5YvAwHIDATg6TfRUtUYMof2d7RAzD8Et5X5UjI6sM7UByh1T0kshJBjVmskuI45DZ6q
ZKv6VV98LV7eZ9kXfI6taIZq3rcdJbMuqXj8N8ziO7mvEydc/ISfaAuuo/Fo7BEnVkf3lmcqzzcE
qwSjCtkxk7uFCILOF/SggXJ5T8gH794JeyjQwD/fGypciCHU42f96UuBIABFsAjF20BMCSgZakQU
fv06GflKA5b+0Or6FrVhijIFuvpSlqfdeb+g/NEhdcCoxXGS3u/4LEsNxRyBrzyw9RlJa/CgRADl
y5p/5Z8wP6qJVDmShedBbYXzYdSLeo6jUHneCzbhr0YA6n4NPzJJwuJA+MGDUqIlXSc6uPZ0D60N
uIMYDy/RQQtfXa9vSgVApXhJN2z7pdWFZl31z0CofDj7uJu42SKmGuCvJTBsGXLnal+HiyMhu6ts
EIco+fyApfFfiXUgc9f65/Dnm/Gr/4lCxZA7JTozTvgNfZYoh/KNQd2AkqBHeZLPp34wbst2CGTc
NdtrmyE8Xnk5vyICDRAycc6T0mo/sw/e8MLZeCdn+2agLNC+A571a35WYRDGwP6WE6S2Vq3Wx+yf
GqjsFcBeeu285kKxbxCLZghsNA4a4qKUY/V3ZiFPYZU7gQdSrwYq37qQJRn8PVC4tUjS0ZWQiEQT
OdNE7VKOjSdbK44/Hm4GInJ7UIgGh4E5ak8V9szNg21qJ7V0OaGsrbzVlpZlcZHHTKo2yWxLaQSf
89iVzC1YROfgWAcsyL/8VxLfZ3YM6yZJMP7yu0D6N9XydosOMZdUfJnYRi2rK/h+i05QWwqjTnSZ
LW4ZnBFgV/4vEMah+XoAzGAeERyIAF7UhimakdC1DxZyOAFIgLLcoX9f7zWP8AWjZ/4IuTp3xs6N
13HY6A+PUjyDmSyWgYeg5rooy+LFl9vtOTaLcasH4Y84Woq12bYYlKjm8EABs3VMksWlGof0AY3q
XryJNo/c71VwZQcmayXkX8Q0kDzjPawIGdQUOfUWO/6fYMdjPJYv28xBD38owskQHpwyaPgjB3LN
xAZ6Iz9MN8xn8BmWJM1aXUV8LhoZOBibjMDrSnEF+t81l5S6APRAaErI1N7RIuyOiDNvzkjqJ0c5
hWNFFNycQmowfkLXYOwYk6kJwAI3aLe+WmzqJeBKgVpJHdgYZKZ9zDQhFdo51ZrO4/Dbc5ByX15g
zC1kEAxKs0Lb4dO9VnUUDrKTT8evym3RTZ3vZrj0KrZH17yTkXIjPZgkav/M+dKTAfF3HeOyXDNb
vmZiKS1HOljbGFVNSTKhjh9qxcgPhEtF+FCfs3u8d+sbHrEZfGSYTDMpnlz32eUr7LqzSQ2gG3n+
pt1RfmRPWDmTKEDu5rNMdZp2ccsyc8TyxNBVwl2CSxk7sFWE54xGeNPkE+utKrVqhoACecfijNLW
rFho+/uVs+tivmpC0m/anFwGTjOCVxP/xI4sM2AlFadzUY7uZWa1o3Hh41zQe/HNYc68NeJcdEN9
8KfdIyyh20TgjPfyHQLFF6PPkWwXhv9Dg7lumk8iBv1oq2udUsReBVxX1O4yP3bIlrT45WjwvWbT
9oiziM3xSjhTiUsLmma6t05IYkeWseN9pQ08TdiQOQLtZj71TL2JMUFWiUz8cTJhDxPeY5ITczSF
5b9g6yRgelRTVFwTC6jMvK/FAd9cyPwUy0BhP3LSFxUc+gJ/sTSa90ksC+jcCovHj2K5InFmdeLa
fY/nekH7EchqmIy2VLNXrQmGRWuzUmzt5fUJdFF/sBTebcioa7/n49YP9Pbhz7auqW5vkFQVgCKf
qrCqfnCB3ujDKrhadsHJq+y2wrz6W8hkZJ0h8xM/b2aFn71Aoqhhn9j5DZDAD66Qf/lrsvpMEWCf
iGz+4E6vF02hMCDxeOcM0Q2Hf+HPRMdj/8nsMyxZTMDNbFeV8BKu46Vvh1voNWx2cX2cZnqkGOu0
3Vtl5vM4nWVfLqwacXuqSmaHRGLVWzM/oobxNTUIrkyQciNzMoR/gKoZiD6Wchdml7zZ1hiIHa3R
ddLIeo9iXB9NrJeVWW2yiIApjZMVZaPa5oSqxzZsToqXnYyxbdpGR9CceO746AjW/yG/ILK4/6jN
TxEt5Pcdk5wF2g9VMsrOQCZ6lmkDqXiJFioFY/pTXd1AoreXUDKNDhiqVjBnvNW8wZLxoJSFBqD3
B/0Ly06/4eSOxRUj8jNgQfHCULO1DQcYVThh4/s4xyAVRfyIHLrCbDyT/a106F3NhRuexVMODjTz
jU7nbRe8wOEU2vHHJ/gTuE0vtvzH+ARoUzRcSMPl7zYiMwFdt7xu4ZPn+79Y/u2KrotxdnIkV5Qe
OzyHzOujbFKzCOACbBuCSgA7RS7FGk3BBZrIFTw9v2DyAhLPXLgev724udFnDrIBag4JD+THXPKh
vSOUdxuGU9HxAUF6HuOkC7W+ymOMw+m+QGnj1jsEStbWyzQNDN/9K5BxY21gKYCztDS8WXnIG9yd
ascjD8luTWY22Wdzp4MA77qezX/4qnog0dhHXDm1E+u0E0OBC7LeIrL1h3HxZVg/+nGcuWVcFRYj
12xZocrq6A8UlXsVttJz2Yaj9BawQ2TGXUTXqI5QJIPXafmpMxSbUqnSmHdAEBaA/U06gPQcmoJS
ygfVnjQ0trcLV5CDFcEGxhXZSD16UzhWDzovUxTqU06j1ovhdpr02KAWBDQ7MKpS+6fKYqEXsWuN
nyc/W94bhjq7J+HNqfgSM0XudD8hLmb1kJRmScTEBMWazOAYOE8c2jDk+5F2TSqVjqXZzUETUd8r
l1fWw+0GJCHkOvFvmmWkNE0nFrXq6X5se/+1XpjEZW1pyK3A0U/R7NTcubqUPU2qXWixqwWegojw
hRTgdFik2J3LRgn9hnjnD+Lp2Sts9aDrmqj1TZFALLXGwA0Zk3LkKu8vzKE4jSY//NuyfVcBoE65
dqTCSYZ8v7y2mKnqQe3KMLT+0NhHDl251pMxaBSksX+hwQKrs8sdsTBr4CLmaMhYw6NxdoGM6mqp
d+HMYAtGJFMlxJo+gOhuSJq824GtkAbDX6b56mMePfQ7lEDZfq8gGhzCR4jbqLtQWKi747Y/Yya2
QEILaIv+KkYvZF1apK3NliUfHTvjbEjEy1UMVRiQogCdLNCRIknQ1tuth/IPBzKyULSqrJSv1T1X
tXG9Aam8ZBhSNO0NFuCy4xFUV/Z/+tWfc3q9EZlURMRmGeDNPdDIeHPSK76nlaHfoQMVDkBwMoDX
t6cSlIRAHofLtnwQ6J3V5tbdUDINI8q8e2yp20HM5vlfTIdDiUTj1v8k4hE7w5LBBvawPr2jDtix
V4lr2NzPFWcTu21wRtDKZ4mbNmVInUkHPml5Q9wbAMiYWyT94cGbQAA25V43WM5bcMzMtvRYCOwL
5usl+9qs1juYRYRu0druFz3+hETvteg1hyZbXMJVlm85zcwo4EmKLB3dBfpEs80wAjjDNR0lRCNq
5e6j41Y0dO9jEv7/q+9Gi6XdJSmYXFwSGBbo2/HRxMTC95/NkeBFsccM4aCFTF2FdJOqkeV3O/WK
byiuEwPh0VSBdcj3JccOyUeYPBkaJm8L4rt3bXLmWmlR5SlQcV8JH5i2mlsQwYgTzHW/JNroV7OK
F2h7oXiL7brOLM5/BhkxH+4NHVEMWDvmi1tkh398uCRLRGJLse5ZqynnN7ez0IaVHPg1vJ9/nNWa
UqyeDN9CK0omZJDfamKOVS7XcJhIfxCkNrZawmStiVuncPrR8o30EjmeZyi34Pn70RUHqSVrl/5q
cu4aB4Z52cm9vH076n1DG/Zc6FS4BiRDGiZqRh2RPg12f7LblToTEF/w74ELRduhM/5HgXipWalH
Xg6G2sPlshuW/LYG89eL3YWDwdnoMCBR/4kovfYyIJmcloFLiYExZwW7e/g5LwyBCCM2FnAfcu5j
ZAMMFLn1eDJxtW5AA8Ll/XCAxdA75LEU3ehUXEcihsO+uKfv53qA1FYAK5fQ4IztEyNUQd6dthIw
3hnqo7CjOiia2XmgnCaqVvdGNw4W/82ys3eLOFLN1LlN94qwQJ7HtX7Sjl/t+5fwWVWDIaZJr6dB
IZzd3eSPCQiOa2C9Prfpk3Mj4FMIJ1pwnbU8691nDn+559sxkLNHi0BC40gBMlnhrLL5bKEJGNhV
PJ60IJAWFBkPcer32J6DKRhePYiwjA3VDvaT0GJ242l0h6XQoFrEttuyI2nKl0CRQMyWd2+ndQfq
gm9GtswVYoN2ivTgiYx2D9APrp4/ZZqpsgfLal0vTeBd4RWQ3/EKTVw8zsUZlUOL3/oHq9fhI485
eym3gCLF0sKLJXeOd7uHtn2j6hVXLmO387jwfCLHGw3Tv59XOwyhdiaesDkGde2YWauZUCbiQsTC
MlNH6mZu+Sg3LII2u6lsukp2WQVRx3dzkN4vYW3Kb36wdL2YCj7uth/F+/e6stmdIXmCVmp1LeAZ
g3zBBcus3n3nsWNy1DegpgbzkE+JmNSVSi7/7YCvShshyq4f9hQYaNu0z5PyHMBiH1PUL4gfAGXH
dH7WEFseGG7T9WB0wXP6QCK7ECyYNioVeZbrzgfdr/zrX3DDsA5XEFekXH/Uyp9Aq5PmQ5JjHjRu
KM71SYxC5cMw9dTRkm6xCaIAm36vhsrj+q0lH/CYgptxMGbHiNEBvfFzwX5V+kU8Ky+PRGqlySxR
JHDGsbTr9RgnZg2jVMMKIbHeXdVvZ6clTtglIW1Qds2UW3ibUHHrKcd+bnH/xHtpunoGaDcBwyRZ
JCobdni8oeLrwanOHL287CbTyiqDuYyNnBS8x2Qkri8jvZqh5FJyZjvPIHKNLeSlIn5ldTsEKR9S
C9lgEN3W72fY8UowYAt5NsAHvwsllZe/duRzjedoMalXuYLaeHiTYnVyg0qMIkcsy9yKXO0OYZlf
4y4ItQVirGtQ8eMLhMIcEvT52HzTdzKplGqCwuapnpG/I7seNjneXP1D1PILh9S6p/0OrAm9EmsA
vdiD0CAtdZxD3TMl9vzK0uC/6mOvTstuqw8pSN4eUxOOvY3YqGLYZl7pEdFJQROpiDj/HH8uiXl3
3Xj9ivyhmvT7wHpWsUUT+vXRjhsIJj6zjqGOagI8FjmJYGLuMa3ifYE517nROD6lpxL/yWYlo1+r
4Fl6E+IChI4qQP1pEa0MZNQXJLJdxzoUHHeJBZWz36PkiRskzXs/dEtvaHJ2njzp/LjOPgIE8mdp
hj6OIZpaDttk6R7vaTyKzUjtkpjXXrQATKhRwzG1T5jrTUqfUxRcSYrWMjeKNB0SGEfvcLWKlfzK
1s/ZkRYkAKrmd5rhLf0AFMx/fbF9xTk1WlD6UfE1IDj/1V2yvMJLHHxiK4Mcjg/sFZGqRe7MSLEh
C0dGivpiH4uO8ptjmpc8pd4IU/8M63CGh2MbKWIWjzthjUCPaymzMHzuP8OpJaCLEvolSeNA6ZmD
I9RwoEuzvXq9wpD/0h1piC9HXxYf/BeDo1hcFQfmTGIQTFRV0bD8id6Q+rulDtRlEdGoGXQo+/jP
WgUWuQKH0PNl2Xwwfeg+T07zwp8HalsNOckeKcqwWq6ht7lp0BXUInJACGEy61Pviz1BUvn/SPGI
46kBzpQeKc4ChudRu0iubrRJa2NhDcyuBw1jBhdv2zni9W5sBhN5OjpEB+dXcy/I8KSE6wsch+um
Jr290Lsuwd8w4vz3K11B20sug21p8RjueWGw13723rPx9sMYVFEHuW1xigcgv3mRiQ6G6hkAFT1u
3rjCHfvB50so150ZhzQPtK1J8fkozydkGhsE32lpL2JBVNlUo2G5ItsIBSmR6ppblYpOmebY5dr8
Hx8kAuqqblpVpO8Swqlze8IoL/oUrZH/dXMZGsIO/tTaFNLRgctmyR7hluItQ4GzHwjytf60BrLM
qAlQ8yzgkO/zk+M8MQQIp/MsoC/cR93GEsFnP0Raq3+40y1j6ZM8AgsI/1zSO40fAXHWMiUGsiVg
m9Ig0TNrgu6++6vCAvv1RT+BQEv/FYJmt3Y31+Ul+8kHh+3YRU25SOSYtFS25PpolrEYWAox5T41
pBjdk07vOE3LDS4S9P2yKuOdKSIaGvRkA3aOVW8EeBJ1FPanfBfDXEQLRvuORxX81NrVKFKyXuVX
cSkNR9Jdj/3JSMNwrysf/Q7Qxl2mL40I4mf8L0PIpKLk4aHuXaJXcDHgbJapfCrrEnD4BwsR1bLF
uGthUUEcAFvDmVhvvky4PAX9TxNaxnxdCSmpDRsMDZmJNsn1KQv3dVeX1kksnqxGmbTmdX/ywNGT
LT1ZkkdIzf7l790kJZrpykc+jI2kFDCsKDFYU16oVqko1sHZOordeaJofohhqOQSRfKxA1XzdSXa
fH2w5HtfKzUENZr7sSw3/RxlPeqAwNmNUdA9S5C97OHZojppqyuYsJiAV/+ZIvq3TMX36gJuQB0U
xY7qqhuJcbsgVgo/jQPJ2XQDO2WqAY8gAAwW675LhE2MrqWvTt8CNqASqA5BETeRFHVSqQCX9Idp
GO91Gr/haon/0SorUR9/C+xG4DyNaAud4Hu0aBIKVfv9xfpntfZi8FvB4hk5cDiLAtxFnE0jIWh0
UO91uUUk/zCKXP2Bo/8PAg/7pT7ceiPV7lMPYWD+SxVWPRlSkrcxKQZoOAxO6+x2wnO/q2Whme+3
Rn9qXdmDvjw3Bb41H0rchNJaoEGwf8PVVtG+nqI+kO4qcHaEtTo57HFm15HPQurYwLByvSK/vBaE
OGp/en3HEz2EGetl6SwPc1rw5GXVpKbHd4zSlK9N0QYE2l/kjOWq7cGsZNOjtj38/xfdnzE7rc+n
gMmHu516gd3wkj3F3C1EYYhvT1Og5ui4SUoVM7EKMqiSJFnsNwVt4rjeDF4Q069xKa3ZIEsZ+pZT
6CssiPso1ci8wEzTZ3BN1iHzizPqi/qDig1IRPSjV8f/meiKP978aNKGR9YA0LPCesOKij/+4q7z
nDd6dorMx4MUYeQ+QNqy1jXg7Y57J5/SKVTFxYQPWeIiaCuw49VQ9rPoExP+ffLcSNUytY+bjr6U
1o+U95QzRZejVP6STBgaqXicmNUzU5mnCtlvVOj/0ufx/033mE26HrAhSLLIMG30WOqY1F44n4Nq
rRF9gG0FmrIZfFUPRlw6YYWXKl7T4jWWIdSMQMfMGloFg6rWQCoxjdKLKJluj23FxownBIJRR5fX
lGIs8mwZBkXzsPwuxpXAKpFm5Wbx2pHDekb78wfeSTkdxqcGfw8b9OshBfINBeVrJuqK/V3az4+e
ZWujFraIpbMCVB8HS2zg1vYQaCE/wVNUgzUCm9vrjgwN6dFgQMncBM1UixzziASg3XE2N3Hhz0Ld
BJSxLUUbZgu2+sKI07nTG3eM/F28hyjM8J5UM98mnivFAmrhNInY86DShJcXQ1+qB0YIIRT2QiXD
Eci9o92qHCvzJPj6vBiZTrC9bW/mw7jUo8+leNvSx2Cxlh+oOXy65iAiIZCiCrVSRX9YJ2z6Fj0l
YGd7ixinO7Ks+WFoh7+UqMkSGh0sIS6dwaiz/I74nsadw39pnJrW2t27YdIW2160gMQlNm0Zi3MH
7AnsNpwXxCf+W2EQWrHasD3swWSlvOWaqLL13bvfGQmA+c2n2QTrm2CMnyFVXAag/tyvzBCxgZGx
PY+2PL91+QyoGKo/hpnyr4TSFs858rQytWEAL3jWBG5dmdP7zdYFelfjaGCe+fck05kxzPpa84nB
XFP45QIpnNlFKoqgdLDPIowefQXZ5Qocm+AYbvajWb3z6mMS+x2M0pYA5JAE9xC7zZPeCXQFR0Pk
Np2l8l8mpgmDMpptYwJ86xFiv1rpEPhXZlJsXr3p1h8OhvY7cMZh2iiLov24GB1aXLuMx++pcrdx
fRtGXzDjW/wEg+PN0FaaKSMInHDnffn2RvXpm/9E4sZht/kuKGeVYok5JoGMB4nvVGuw/ZC0ipWG
xMi++Zr/Gke0gxB6nGKplL8SK3r5V7/9nwI7bwa7B83aKjtBVkqS580qTAUSCTQsFt3QOO6NxJVh
cjGKtis84p2sQThD6q7nIjmno08cResswaMaBqdkZpPERzMMmORtFscpHAnPBM6+YaNotqlJ5VMk
7R8K77wrcn5I29CcCs54+aMurSwlm4pkKoxRXcdwgx026OLQIU5Q8QlDpIjvX0F2W0zpYjvuRU8m
rfUkwLSy6wvbrk8omPdlk5FQqVl7AextMftf2O+FCuew4C8lrdrNXBhlcBVIDf0bEiBxQO/iriDy
d5KRpZWueh1qIgPHbBBaYnCVbr2t45yl51SvLa8gbZvE2iya+MjasaZFJUSYs80Gl4NR33HmevuM
ldEeZQ+8jJFg1oiDyxmuNjyTGQpXx6RUKuzZB7qg6kRCXlq5KKnFSqt/72xIYukw9HdmzFp4tRBM
ZX4z+FsK2sB8X7rprCaaq+sukZEhz4OJlfo7lgzEs7W8h83cH6GWgEVL4rO4z5OT7AlHxIGm3tO8
qWfDhre0NEZ01tK4rqZ6SomhTy8yxKEPCyNr5G9bqkM8XrPP5r4/NDRkDbyUT+WF9xYQksdVmZGG
xBQYaNNBSP5ZOVMyUedaKJHDzVE6/I0lPKa7MfMVdueri5hF6WAqo05iwRmga+zsTWyCn0htsclT
g0mihWQht7YI8NKgCZUK311wIbxjgj0bJ9AyvediNHgA2bohmHtLoq3ohmegxpeb8woZujFuiU+t
OX7dS4j/lxVtbxksb48IsZ3oBx7yPjW+0qWXr62IDlk6S7IL9YwiA9d+0zC1DYHS8EysKCKn7Gnk
wdq8YXtZYr//4ZMAhDV2ld94dIxhJbiaJnqoZkUpSIefLBuue8EO+NHQwaPu5DzTX8E6RPcR1I73
7IpjI1mRmTvbXypLFumAk6GTioHS4DZIXBhwDD5whkgVSdg+9xeZbAY2AaSyT1Q8lmCp7VaBrMz3
L8mYBs2e5Anax2eKPXh6qkuIutumXs2jmyuFzseU28KCUVhDEp9iuzaF6LI0G94SYxR55kKne/+q
vwQ/FbgLIyhN7Nd8UIAQq0O4epX+vOFh56N9HS4kwMSlRNzHPwMybWc9/p/G8D5/fOHG/WOrK1GI
bHgs4kvkUbQSDC4jaduTloaBdhTkL+4S6G1xy5U7Yu85dFNTbtE589Z8iVwGOohj3ryxBw4dGyz7
Fv6dV9BXbmaJ43BIksEa6V0jo9CiqLnE76u0Dc70nUPPxTjEGlJbkoUJ/EjZpOscRfznclUyeLwU
6yCWzWvptzyST4gHgnBOSsLztxb2AxDJXvqNsIDieBkLzMCMEOuNnODMgbQQlAaCP9NkWF3qzWCH
9bwYp+ajDFrGNOiUMMzVaQHiF2jxO6om7LGuwmh+biVEyznd2azl19/gYLKlLyzwEjo0ErTNgShn
9/iTkUR3KbreGtNC+L2mixKMgnaFd8yiRVk9j8sqevRea1zaHDmzqqPzhEDlMx7R722ORCWgR8Qv
0vIyj2prNDLLIytUOvLWaY7xrMfZwinpEdjgn0enmG6AhF9djqSJ9sbEGjGatjNkYMqJRNJa1tCJ
klmyqw2JwAcKlNQ8zh5HYlSxKRBHBOkxJOxQw7/rOJwwy/uwK/qBVFn9lMgvZftncTZg6soYE9IU
sQ5fEMde9EmFrKrwVCR38vZTgLX869dt4hjkpVpbeoQWDmUddnIIs4+B2Jq6SCaeyoO1iCNwM1Du
ydD+v9FW+i1VL1lMdq8qIhziWX7kQbnVWF0DfXQJUCYMW5EnEkNYLjKzpChVzXon3cxIdFEptBj3
7tES0xP/GpqHnrNqJyFVUW3qxDjJCuREQDkS1+lRtZnKMhVm3QTkX1h7uZoIhmw8KIQnVi1K+Vae
hfySJ4NXlzF5fJAkTn5kGN6erO9J8bor2ldRCi8gdvXmsJmrBIz/ycce+2S8zkH0GzsHtbNz4yfv
zo25L9Ilr7MIVUC3vQmHq8clN7LPHNjdYSFgjw+ia0wUcrqpaX2T6scvRs4xaAp6DIYBH5eCWyRd
XLCfQ1QxTOvzI/nYn7odjhYqfLMq/RKZdirwhZYMHkrcDnk7UvuAjxJGtUMC9EY/scg+aCL638SW
aCNCL6uanRi/FgB/Y3M4fcWuDLeEMPCQCIGb3hfq3MNX0me0C+3loMnf6Q0QGgMD89kkAh4aoL+N
U0laGzWjnlHd01vq6bVfb9hYyFtnqZ7mc+8NQ3ngZTlpfX/u9s5TUrx/9IIUey46wAtwl1CHcUty
ZoFUo2fDsXdoDkuIqfIAA2tuLCfpA1ZdzChQLFpCVWOg/KhyLFvHpnm0F1Q6HJ3qJIdgUbOlBNMY
HJAFKmfVaV7Q0WIWYZauMe3zsNUMJyY67aUJdaRWzXnp6tX0+XSocL1tLvhtWeYJzxQmY/jAA6K2
i1WxQgsMdRhwfBZviAUXcnUpkNRP3rJXe9lacKnmpbTBbrQeZznQgPPqdlXrV/1H5M0tvQcsJhHd
d3KQsp3FX2yjUKNdV/Pe4m82ot07vufwUbYxCp1dRlcAY/xtxmXCoxjtWRC0kmD4NiBX0c85UYeX
nrdd3MaiYOme+w4dovMau8i+CNZ2aRnrLUD9kH0lGuKhVWiSUbD0FgBH0vZCLIOwPTAYAQTtVikE
GBIhLqmYYVOqB9wbjFQBWYZfVzJ6PtEA3WkNrDPkBTglMPC714Znn19gNgL/fOITBXjhe5cLKuwB
eilWC/mkThJ2aQczin3hkcXZvCtPnkhmyzNZI//H8fPqsEoYUGHhEaZJkvRvF9c1k6kBC03E+XdL
iMCnzV1tj/ypN00+VorCvy/ORlLPy2zU59RY3OL17gTiqD6X5r02Nn3NMd6ZxBpoSmtzkzg6XabU
XVianaK7lai3xCvspAJdXoSuOwdFkngGfOeb9MYlk7KkshNmcR1RAmfSB+ZizwqIXYBECO9hHuPf
2K/6LQmPValGpHPg1yokmoDHCBEcRjwOmznNN0kREH9g5O31GJwIwX9V4829JEpV+hA7SEOT6kC6
1Qgqc7cVZw6io2ICUfP++OXpv99GsuqHJwtxGDVb/13qk6nbMj1ICiSP5s77t/eWwZAFFLttDYdn
Lo0R3TlhtWrNFNazoEGHrc/Q9gBJ9gIm5y63m+DzK09dtvzpq6NeWWHabPuby81Q50HwiBxkjZMW
OVCTal7auxFyfzBGPhp90wkH8Kt6O69J2+mdRxjNV9m2H3TUxgOB8UqGcZz6WxIBLo7DGzca7fJx
/bQbIZjTO+f/3LZrLS4LgxAEDUkuNdQEnkZHaZqM+PCC/lC1UXsIolC7FtaIBxJG7Va7H3To/s2G
bcFCMLH4ruZiOZn2hUmjRluteVAhCI/gP5zer3NAgZ/+jw+LqdM5/z4795LM47eADyCrEIDaRfA/
qQLsDoNzgE4yt1Jff09DBb5QnIN5oKeSX07o/ZnwNuG8jQKP0IJglaJNs7qNnxZgXmpuPkBhAWe3
UX8C+pgSHlTmzxXA5/co3oaGQy2cWqQmWd9xO0OfRsXDz+owUBQmCmGySHXpQJfny6oMsm+LnvlX
JajhDPtx1N8aGFqMVHrboIzAakdQ+Ya+dXP1BYH3Lt9u6CUWbM7tEzvzbVcVns9klTcHMthA+0oz
FgfFSujSLECtnSYPXZGclXuZ0MNctfyb1N/NKQGpyD/u1xGA3vPM5zraGXIB1jwzPtdDJhxiwaqd
YHlSVZroVGs4BJqkcVAhR6sGcvDC3wPR4cmGCZY3HH4LR6gYQkxiieV1Ch/XjBgmkS5UPWHggfTj
dxWt5cY6pppfQp/nXMKi4uKFMezWuelyGcgqf9KA9VIWJQssMgBZ2NPajY1XyEk1ATXkDwBQ+Y5k
nxM888TC3jj3ZvbFimzdvMsP4oJNrcPMvfIH4djbQZg7HzIdFmxBGSqYspG4+rZk1SNpl4GstgjR
ScPWNBcJJ1WYQnMQ7elA/YCrGQphADdj2UPEfOZhKvK8mjvJBUCQTV/ULoJGH8UzvQ+nj+LTORmA
wYk1lZXER1OBQ2F1MrqZU3G/XWCy6W0S3Hlb4/Y96/IKU4HsanfBaIt6Wn7Y1CB2RNBsfMn+wt7o
+uJTiSTRILvZN2GG6uWjb771+DflrDylkIeZ9Qsxy1ODZilXqT8NAXqmyHyE5Jwofh+rQ/qvkm78
sCFiEEXfulGY1/DC0wB+CGWYDVJBz/qB3H0mnmDUvyAaojfbemkOo6mHXBq5OKHTqfYGZgbyX6p7
VEFyO1v+g2BeFtGOi/TjDlozkRlBYf8DIFF6lFb+M101jL5LLSXiD3runJbuaMWZWVK9Z3De95FP
0ma7zkAxUYxL/Wn6ZDxE7LyTbFhzBwOpwLEvSE15fO40vxKrsyZAW7tkVhNNpBVnIHTk74fMDInk
4cLHOig/JFZhdrCbRVhAl1GfdqLGug0V2Vl3fBr+Scm+zWl0/T9RhciZR3JRJXyQspSiLs1f8r3s
ijADYf95JJ7HdKsV+TU79o01D0JLe7TkO5VHoOTSG41wI3hA1wJtPgCGTWWVEo6TdW6kjuITrJCQ
mKmDMZYD9E0ncKURsHpq5L3t4DROq4uPl05M+7GcfQq9LGyfi79qFu5TfVRkv3np+Q27571kunRU
ND8UBtRn2I6aTdvZJBvNlE3EtMa2GvymracPruwuDD27t5Xuim2gfcEoqAGCJoZCNQlT5eobAt18
5MqkewRp+A/+ubWVuAaBpjc9g3Ma/8bjjjfNLf3Crxe7g7krkcdpGKlAHT1ZpZ6b+gkLo094K37S
EYVwYdJg+rOQrjXp0vWAXoB5UJPOwMc2S7+kCtTDv0cDCoFMFP50tYf1pRsQCXWXNokR9IgzLeYd
d0YSoikrdZlJALQHy/MlCt86VJlhyUS9YjC1NYdpZK3SSMrYua1tI+CAAEtfdxjdXhxNcW6SarnQ
ktTmH0zGv6phpN5tuWbJRsFHVFKI41aDXudGy63wM4LxYXFWMKD64gZp4HdrynAwySUxj5ZVagcH
PtyiLU/55thjMFf6AU9j32kyxEjoy9lI1ZvdvHYdQrI7SpiO9gRAdqU7RueUyt7DOidjv//BjTWL
JTwUrSZoFrjQY1w69FX/340e57sBLmyCHLdeKPCPLfKuNO1usCX24e4MyJ5QwF2qCjEcyhLwKDdJ
P8OX1q1GKh3FqwFAVOWPEXu4Freu2duFPB6EDmAjaKHieRZYmJuyo252cjUVL1gsXDuDu49Cx4MD
cbcUgNS19TkCjLBTpjJBowOQjFXEfTvvHIhf2hY+IvFgPYHLi9V2STmYw3mFK9MXztSK/MxsjQZy
IJzQXV6GPrVq7Ubi9ofD3soghBM8YJpT2zOVlrTtNPONuKHEuAH3Imy5xPoLYK4tfQSmhhk1XfKJ
EAmJeZZNH7wYrTgMAs3GXk/JLNxOqy06HXXPsm/CB+bCQM/NLlDCvFMVyMirnLKzc17liBPYtruM
muEaDyWQkzpzYGhy/oxonY8gqZOhfyqyVEeU2X7FXV8HvLT49LgooWhc7cznKSoCFXhItl7m+Vns
yGSCG7I7ELHTPklFocEGa5l7EAgysq/tNK7Cwtjst6ZbwKYFdJRtll2UTgTDZ+Pw/YIKdkwKXNF3
EVVjVKUqGq0sVJbpSJgAvwSl9cC8lbjUAKY5xooTJLz14Mu7yDwGoFTWW6dsEFdbx+pb9ndtNWp3
9IGwwL4z64idHSwUEyoBe/B3D+tCLQRR/umtq9LXuI6PybRgtL5Dv2Qxjj0jmoVLegHuaflkZrHM
F4SSdRSYuO1/66VnhIUDZpI4nmFsH8psuac3M7fkLBBVu5mTNwXKFma3Uwgdk3h/j2iPT1Fh4l2k
dN87W+1MpkA5rOsoXWwaxVoDtLQH/DLvS+qKaZG2Oyanm8GrxMun17jfkBuJNkftY8T+ZpRI5nZf
mg4JgZyFZx7GPI3zhmDWinJOo0JjROT+yeny7cYlOWIMmcnOLMagWPk2u/PJxvsqf548Z/gHQ3bq
hsP+u95kI80Rf1i+ZuNSfzDGM7mqRzXzAbmIfnZV2ZWq5ac3XPhpirOrEjP9zYGTVgI/sAH+Erem
FQYph6M270TGnqRIprS1+3fPrZQGXjlB5wVTYiNjSrM2om48bx8T/Cx021gdhLqYSg/+A3eTIvht
sGpzl5S3K3at3+g45cgo9x0G5Vv0rUBx/wEcwoOFbc3WZv/VYrJlJO6gPGQz4lawQYSE3VuZGUWm
/ujx32tyGrBDNZbVwrLLiHQKjQeyEeispw1Ms1CZXVxR88oSKiG6Ac1TBjR7JqXY2i2WngaMfLAb
/KzPhfoJGO28zuK/OLRT7BI1MwaWPQJ+8usYEq7/qPgJDLjFYBKA7XNDvQV99HojsniuHtPffkMS
O6lnHHdqrelWHy8gW0XQ3JiXTGo8SF2pcSnUxc/77bwVBGbVdn/aUJMn+kY99rg9ivFfeVKVcwSx
0Y9qWuivjQiNrEOUyJG7++fv4XiLZZmXgnWpwiJYrK7q77csu8pZz4fv6Ft1vaJsodVPvjBUjs8s
Wo/L9AwPJ6qLJ8JmD7Igch27nEcfnmzX8IKlUBbt60F/En7M5BU0p3SONXCXxYvjEryfNrxfPDVL
AMDv2QFYP4Tb8F5Ptvl3nleyQOkUXOfNpywpUIDvv4mrUzSirgeiel1hAPgodyBfHB+8bKh31Yax
wZjW+vOfDeqTmFbo5tvaBym92MrhTjEKu3ARXVaDJHXfL8dS07eDLwJXvH/ZonRy/tRIV+TeOsJd
+i6d8/T2O1dduxMCnTvKe3IgYjd1H5uzrftxBeHlSPOKEtCbB/BTNzqhrHSQJS3ICpsS8cuQ4fDP
UV9kID/IvN7acpBX5lTGC1vPb8bIukhHDsjU9jiEVZkR7///pR/nFxbmmc+ksi/y8zFhhZB3GyVU
o8Q5kJz2+NFVvtB4zi4r8UEkjtr7oMGwsfWQN4HeLQ/B3gnQpiD0jMoli0r5mBm7+IiRW3RZpz2f
22AucxLG8deCh90svG8XSI1LQBPfcUndbB1BjDF9mRlbJXgIyi6CS6g2fBrY7dYeVB/LW0k/N1qV
yio/5dBXhXZ/fh9OIKmFR5bV80HggrmlmNx94ZnkGSww4M0Pj24lgRe5fW8VzLN6SDXpFT94z07+
GNoWxE4DI9FsD3RI7bY6cUxVfFakTYjU8pQtWTefvJAs9aUOzfvV3BrwxeouKGjA5aL1g4SzMLXB
MGMPrh7gA3siqFNoyhYpDERR+tkUS8HuEapBsPUbUZe4HseVfidnAFP+nu0Hg7pUUq6Exr4w0EUL
a5DrhmeerB02cjw6opSQgvkspi0wgf85Ep6SYNajDUeY4b1dyzMIaTE9Bm+ORq+ire3LG2Vf8S+9
xRFdHL22j6WE3mEPE5YaiW9NjN77hk3Qjq0zaN+BBIukHUanrJbzyMrUB9H2zZGtE+qNoB704tY9
UMki7WRl6NNiR9q0koIKeofFawXZuOPhna/sz/Vm7oEacdZ1LrDhgekI6UY4AZUoS8Fnnkstkh4k
FULypDBTMvvIV6ychdUx1QHkzWb0T9k494YESRCVXHMovPlnWyqk4YIjVwdDHt73pcrBqpiMGYHL
m6A8dJ2Eg5mNPMLrQ8p5HLmRfdBdFiOp3V2Eege+e7Ife6Ush3D+GGVrMqSIzO87DoaJ/jioMsVZ
tCnrnIQMr76hAOHrc9oofXqGmeWS/c03FUguB5nvAkoeo3KpomtD9Slx4VhESJqCOkAW7IJ+82Qt
ysYs5gfpCERZFBIsRg0qSOpGcJmO967x2EmUGH1n81USfeUXr525g8TkvxEPEe/T1W0VubkwcJkj
wnsGEkH+52e7SZ+eZgaEILOSoRRJtYE0qOyHrM7iRAYFo19uDu7vaymOkJVcLqsprq+4tiqsXJ+x
z3PwRudKfe/qxm3aR0jzv29kqrOGSiEvz/OhbhLOKs2mGTjiMacv7r36LzJFcHQKbVwoKe5x2j5a
tcQEkEwkmmcq23ltK5gn3QVlc/kosBEx88il64tJv1YIS94hP5j7nCtxPEk/Zm9H8ObdPNQ9m8+t
TtyhXnzl564MW6SCDMTKFeKC2/ow5/cLdEW7eNCOHt6834YuZOWLJJERoyh/swn8s43iBficHCw+
+vPlekM4Rmj8XEMbBl57+CXQ4Q2JjUM4Ji16C0uwCGkuKc11QgJsqRDh9ykEyiUFxX65RoBpYxZe
HbieCIjG1uFwtDtuU7TmNVHMmBTXkkS/yv8uDKvfHjJlFO2ZpqsBGVxV8Q75Vt9yRGI7C7RQEV60
2rjnSaglUcweqWnBAw+IXZmyVxQiqrLMUpbvVKD7AlK/veF7g0VOfoVe6o4CXw/NXWPhAE2zjbwY
IiTmnpfSw2FBE7FiYH50qvkVAyt6T+xlbjnDYqVpbD6vA4ZzjR6gsIwVhEALb1uY9u6fhm9pJ452
bHcxKvRLg1qfujKkPpSnQC1THDPZsvi5QRZsk4t7/tDjx8naOMVzDrFof6L//HwHyVzJZTxCLm5f
oemwZofMk9ogS/AKZwPb3/Cshuy37FzWu0RwzMmtTpkN/57ijgBw41tRAIkaFUAzOUSj0+wIjpUu
s8H/jpJjWSSw6Gu2rm9NbbiACWws6JCI+FlDJS0hYIf8t0JIrq6GS/Vvkt7DwidKZoqCyS+k7WJh
vMfhKVgILz5W5o5/owvTtrOtGUpG9HmtYb5S6BeiwtG043HEOHNVsjJt3AGZHhKi8T20HEx0Do4I
RGKx4K9djdSKk1+u7P2fH1RZb9rJJrzP/2AOXfOm5V/z6FjTqZLSNsxgMUqxwmINTShGcS4tmkyF
B1E9bdeXbzInHe2mNgZ96+loLu5zna/j80DY0ksuzA/Gt08waXFKc1iibqWPUo7onHuq0Xx1PLME
yFdJP+i8ZaORAHxFsi+NLBX9u5jPxUGrcQrLB1pKLjtLIeJeLNcOUr7ZFriAHNghbDKSpPp2v8vq
z9hgGMowWRUN9F49r+UN9xDA8YajB9NvxPN6qs3ILMdnLxFKbO5sMnvD6MkNJv/DqcNFjMh46+lm
LP+BhW3Daw8L4RE7VD14w/+2zQpvQiS9Z8IW9N6F5TzDIwmHMdZBi+t/9Syfbi2gZLlFdjyVbDWT
NcXp3cnO4ZjlatMM2smTJFzhBlU74iX5/5Nl/Go52WmO12ub9CnTShzHMu5gMrz4TREY9yLSp4g1
zjW9Zpzg0iYBt0f+FGv6lbGCXmkc7XjKdv/M+v8hSH0jyYi86H3M8eMbJVnOd9e/bG9cplQ9u46Z
Y+bjjFOdSKryYC8vMj5wydc9ccpz6w5KnYRZGGhkor2C1FB7/JP/2F5UapppEynDoXkWnCKKa3H/
XfHi8S0YyrzyFrNPnDa5/QYPy2yT6N61DdznuTm8qg2JiYoDZrwkgQXqDWYrVSVbuDHSJ5sY2dzU
OkfWfsevYIt+KHammMwuWQgtVvUI0V6FuUqX+vjbtuqkl8atEbh8d9XZdjhJJMSjcJGDv0mmw0Sb
cCzglKcMxUO+adK46qsoZ8XdRvNV9dMH3kcwwl944ONe+snzfJ/Eo3RFgIcXxf4V/ei1wLjmP3Ca
LO1+Qz3AZtU4spd38R3JgKMIgBujYh7RdwVi9TcFzko2y43hvlTEObJjgxKuf5Ea/ZhJzvXtrkPo
0ybUFXda379k6+MIemv89pj4CE4Q6pySwVbhG2JL6u5IRU0AI0oqsDmbTJnW+MYmgfGzsiMCnSvJ
dU9OhgIAKNgaWGJy3vzFlPtUF8xdDMCN7I+J63r0tSNddY6bQnz3VDg/X2v9GD6mBRG8g26A189+
mHOI4kYuzmVyVql4BlqYan2ZzClYsJq0PMFF10wgJ5iHF4c8en4NVUOvx0F+oK6ARlLrjYy/NnCc
a/IkShV3wku0tq1DAZxdXF3/SDLxQMlfinn3m5VMv8qMYGm1eLA9zZ9CjfD7KsvUOJ568RQ6Wp1V
XZfHqoe6a/gbl4xRcluaZS+gNUzIhaAipSvyO/+5Tx0oP9Il5Coh7Hr+4k/XlfQqCTphrTBzwezX
2h6xtlDOEVOoObfny9ZhFreuc9SFyuFoabOpRX44C6az99GPw/aRifrR5HGXa1nvafEPc6nvZDWh
FxGAX8U9WufpKaErv2b536SnruuwySoCsz5wh95agntRXTO044ZjqPap5MvSShJbV7TT3VolUQ9s
u4+l7z/t1iUFz/GO+FoUBIb08MtRDVD8FE49lXML4zZbwxiI5ry8m1hqafmkwk0KIKuv6ZgTGok+
3VaPOrERDfHOAWC8GfJY1WxyG113sjlQbre924I05dY2oqd7bkddTD7xQI4GxSOEpHVqaRJjkofq
pYLuzgDcw9BEm8gpZfieP76HT4DWqiVT3DRxcE1Pf71evv9v9JpsTFkQWUDj435BK9M4tA5CpwpY
SNLcBL6kz9kBRq2cgr1zWqr7+XPK1HLeTX3aT0Sw/mznf/8mcgE80ETdguH7PmB+jry9YGcCfYMT
oul+IUoVEyAuZq2vamnO8ClK5XWwfwNYEhwRoSYNrlN8tTjNNi1q4az1+fSu9C6HHcWUv8BEp3NJ
sgW7oETdEXSVB+5Tju5z06Ql71J+/4vycUSPja9HpByFBaRdYMZsS862hnX2jsxWp1ZhBn29XhDJ
71b11ak+me1C/8jEv0mukCPmzrMBJbnxcFBMeaK2fwJ84xDJzK9GL9Yv6NHXO1c5uNW9PI8Azpyu
ulotp3tfeeXRj8ZNC18VFse3H2bHVOz1CaaG5wjjwpjnbhT322RKmLNH0AH/sNKHgYYlgtQ8wiWK
iU82mk3h3QwsPfhr7CsuRT7rFiBkv55ElbCfoYvrPAMFELDdOHnnd8r6X/6nFj8jX/szhU9TRljs
GSicZK4vFio3DXcYp9AdZbHcYw6E0+Yclt00gbZHdwIxprcZikh3NS2RZSv6c9FHdjwgu1exkIU3
AXaFXPMQdt1oPe+SKt9VMr9LmNX6IfhVg5hDZJbWYrzDqnQesGRMtDKi5YrW9fIbt4YNNww0s6fZ
PqKsKUjokJ4uFza58rPLe+I2wxVGY0ZtXtbIOehCiJgJMBXnrGkGLQ738AV0aoX3w8xgFtNL2g3l
ES8IpaJwiS2tOqTq0IIFlel5Fs/0tqiD3lWxCfRwz75c1IJoVPb2awunsgChuZc8H7FjoMdwyVsx
JMDbFnRWiVyjMdp/MhiirqJaZkcHZNF8uiR8Sw8HR8DR3ls9FzyKs+/skjgam+w/GBrygPzL2nFi
xPEI5WTZnJ6dRIgzTRQaKYUnfpDwpJboSIHQCiHZb4o2OmjCydUnVM9i/whm1kZF7EcK/JN4fKTz
v8Ld9G+fo9kkVPYHVIKVe059enVhrnIGf1ci0Wx3gKEj64flt/v5YvSSh/qUPebeFsCIulsb0+2h
SiyGnSmfMh2S6QJgCgbX9y/LBdTNa4M8tLTj45xrmw/blfHJCt5vUQLA7h8BkKD4LcNLEYWdGuNV
ahVhYhLzgTYWmATOEn0OkS87/WBiseG+b0xyey+ZqtusDkY0yxg8QjvNxv5TvV3lhgHKt1ZqSmBf
aDFH9jDlGqbqMhyRXQ38+dLT7E9ITJK2XwjeoY6x+dVsmVK60iSGDRrAEYC19dLlb08j9+2aNl1x
jePCW3azG9Qhc5k+iUJya9BaNjHIlnHAfzuESweZN112oRgw2TTroGMJZi/64S1UoREKRNKTsBQD
ypiIFmvnajPCWpOM+dF+OhskXIufWF/ePqJWsE/6T/TAYCbGJGdDfov7KTXBsQ6X+xD9nVQM591w
KL4B67mnqopMzSCApBMO9A4Dm8VSSosluDMU0m4ky/VhReDVlGIU5hDNewyLe/KAHV5thVdPexzI
1OeYaiQAu0TMHJbUqUxomwl3aN1KZxBAEhuCcEEhiOpwnc0OgVfA5tbyXIUEqqT3QaEpS3lMjZCh
tRX0CyP2ukVd1Ole7XJgT6mBIuUbL/OW5IfXX9HLCnVNG0DM7tE/kTzeW+hqY7Ruk9CUSUYaDiM3
7NnXpr5xkglZYqP+Xc23+1fhiaI16pnL4QeLUKSTO+l4Vc8Yp7XbNH4ZE27Y7poC/7neSjAFBxp7
2IugEpmynJDVE7WQJ+NnnHhyLK7bv3PVUhVpbXqwdwtJ3c5RqcfK+l3lGWsWwmPQFexHFwvZDW5O
TQgQAUBd22WPhiLSdC5bTNrhl+uxDxTkAsZIP4c3tOwfE/zMirxD16aWXKQwCdzeV4nK0p4I1DPt
HxZEIDTGeL8OR5G4xlnMRrdKHX6MSLk0D6Yb2FvhQS7+f2OzEExcajdr/SDjP2NF+vlOPkfagWBq
twg77Iv+3lQg1XKqL7oiU1fXshRuc/Kc5ETfu8PqKLjEKZS2Sj4OqUFDlQE0oQQQiGluXOLhvRLB
D3QJC3kmSL0Zuvy2Wlv0k/awtMnmGkB2g8/tDUudUO3emCqjK8qZ6goFPWn3ZiVv1ztNzFOfEO8V
GiJ2xHM1Aa7BHG/3GDCxOgZaWAf/gl+kYhw7c7mEdT/VDvMVc0diZnXfCd8Tj+OAjlK6uAoc3Ggj
4NJWnwCHyyk1G/LVSuJHkIs8CHOqxaT9TB/NO7N78mP2rxwN8zskCApt4A0CJ4Jt3jcImjS6Rb40
5AkBqQN8T1S7NnAo25YfthDvdyawDd5AMTteHfOUtGl63oVzLEHcNbg+BK8LYgI0pW3RnU6eT7kW
eUU36o2PuzpUc9QZmQvXb/2SuglSlqMFbuATQPtacxq+zy8yLn4KIlBa913tg91EbV+d8qwuhjDx
n73BFvVWvljfKdJARFqyWs6m18yazZb/Az1AdkXoOsJ3zb5+0Xo0LYRlspove6seqqVW9Md/t4Cn
6W3HdVBbVHooItiO/rOsuZgkH/Nm461ILYNwSPmqk542oz0z4Tge54YQo2Gu/DleF+/QTyviASEt
Fxnn8XzZYK88+k/5cFR32Iwf5+HbObXr9isrD1z517IoPfntTBr8B39046bJi0JhJJj5qh6eWCNM
FweQd8vPorlFj/8IMucYj/FX7Zolpo2rHa94Y4W9Fm7lutH8wQS7/oC0b6/mDNgU3Ejt1/SSI/Ka
T4NqDMiWkXMMHPN6jjESsP3kjkRrVWfURT+mLUg0nNEAgB9AIp/sGUSWkj3YJpeDoPlqPrP/lGTe
0qViJc81Indza8HcIpZWs8amnSR/+8szZRlXPCbVuWHD8ZQzbW3r6wzIPJuu8H0N6kfBbw6C2O0x
KC8Zo4XySJownBYYgYg1IOr+m/62at0dsBmq524dvof5vaFnRQAG4P50xpUocnibVMDBEal9Q/LZ
fTqvSdC+Brm9xo3wczH3dVdF5wAgiq0hmYPSBfXTp7irYP3gAW63eUvRBcfeEIlScHff8Sivn8gK
G94Xm/qhbGlCZ5RsAeGNVyGA1niNsimtJTeUiSZY3S024/r2azpfJWfc3PTm0oK3cIjuzIHgcAxv
nfinXYUIi8gsv8zCytQihW14GwfalTdCggoeyELTFMw6o4aRuHrU3iW+zf2HSs+qsBhQhX/iXMKg
UACcHdLIao59gQHFWQyKo6qk8l7VsXwnxwXZgQiPjNDbOhfXWkwCC/6rOngEXzr/IWaaE4afgHAo
VmjRvWnqQ+fJHEDGSX8py5FzJ6SDKl7lKPW9CTsvR6zk847bv7p0y0Du1KBHcFOhbkSVzTaQhmUN
dYVSx8OO4tp/VnTE34U3Re4rD/UuT9KsFT4CMcGEzR0lqFfrgCn7tNbwnXSexpI2lvK1H2LGY7aj
e2ISiqWfZ6CIlHE5g+nmfvQfPqhdl+HlstCrlRIqPO7EDglfZFhS7dl2i3gs3JpMZkziNoBPJnZ7
fw27fzzITwyRBF1or5+8Feb9q6PplrT4A5fEFQL7jeTAu5kPEDSO4119fRZvp1xVXUMqyduoyLMs
5+dkij7KMqZ9uu1QxukVs4A09kas7AMpoQDsT4T1XV2g1eFEMlVjOV1y8HJ2jOeE7brhLD2nv+Oa
GIqsc4a/sljI0Jd+85IthZAVsBSYvvpySyV2FscpANFRyrJqDsBBuapOEG7hlcaB115b2CTc+mPH
OttkSXL/63lQGjWrhpDeM1qmM+isQ+xhyH2BpFtJrGb0VrjYH6/M64cJ2hcI+JogvfJhXCilufE0
GKUcKJzHCObUDqywtALThvyI9yxsGnS9HbwqGU/hnjujax1Lru4tOCyHM50W5YsNGCOTt6tcTxaI
mhloIdNaG/zCTIcJ9z/xLXsCP88PGmFEfAEOBg7AAD8CMDwQVYkgRZQYak7Smo0x09BewRxEi2y/
GG7bn6RsFrkCm4y3Mej+TgCfEhpKttoiRJW3I6rXFuynQx1V3SlIvm5UJy8YD1IW5YPAy7RRi96S
LMYBubmFb8kfQiA5RMesWmGL6TkypK/2wxdW1X3nF1J0aYeWvub9Syt4NlVihq1Yi8bj38qwumij
nBBAwBCsGg4RceN/AFMJY10Xx/yiGRNYBvLDtLXedRlWtzzk6l9izPeo2kPAQYLQbrv8xxTQbbUv
zvY8b9b1EoXje2mjHUrqQ4mSBPfrUS3/g7RNhmW7V/mWSGCdwcqwwdOdd9ZoYfMLfAiE+7BIZs8+
/RmI5D29RLOoYRWJ9UD2fh77Qb35zuihIK+8V2/zmpQ075HK2xuUF5JxIrsXP6wcYUs5ulQpc3Ao
vSZPWP6BCVzKMJpYT0bJquMWNy5sRUZrT2DfdYESLZc2dsmo65OS7IHphFb0GP1ftw0IkWm2EdZ+
bs4aWZbVwSscPgBDsD4NWLbwFZ4KllMrLnv8fgtgyUsuaqMLi4mvF0c6dSbSssmpZanDmFi74IXG
kLlgMuZAfO7rdTkueQIpzBoB31o3M/7WX8emzMDyDrDYWHER89Q6qj0k8D+88YO073HENZoDsqxs
8MYPTqF0lNvP8yHLQSp/LPJ1aKLaW4RPgnq00GozIKHea8C5gbs7AkxhnTJp7EElQo5yP6fhalxH
owiH+nrf865geWSTWjVqNc/B4PXYBpI+eDR2Hd3paB9hu3kMwtLBdT0UZ+48NSbUOR8QRtKcdpj7
7Tuq3XTrVvL3iXfcabSWRLeU/ZTbXJbhkOvZ3r+jz5CSj9ixkHX0y+AtZ2jFUY5LZ6pVy+e5oFK9
VdQCj6c7+/uxM6sIto7DjbAHOsb4UwgYI8n0Pk7TlxMGDtMriZZ1uB2BkRKTvtUgxPA4FlOSlGu8
IOGBy61AELoS/rf7+giqVLC0k7oZ3MIcqO/2cDAKtLikc8NiPaxr2+D4K2gxab62K+wlfc46zRep
jbcbFmNYrqV735sJcF98J85MmI4wUwGD9o3Wvc6kwblJwaAh9oY2LNFXixAenPKyIY375+k05z4v
5UO8kjX5AcK0FBfgDEjmhgRPPR49t+q57GbSdWaCNCXUdiCZtfv5KZD6u/k+krqjDMSxjfHx+PxT
8Tb2WgJHneweDVy8xw53JRnTM7dgcBaVVsAqVpjF1XktVtsQMWW640OdFpG5qm7d7b1vHwsr0yTh
xieT/F6yAyxfoOAc5zv0dl6+iOTEWNNJZhMl0NFKvda7/d4HyuMuwYmJavxgZK8n1hOITtAx8Fv7
O1owzYsIwM9jm3DM3CEObPeS76BryPSGb5k9SMa5AUCvKqmQ7O4/LPUlMWcrixG+Uy0v8n1SCF8Q
PN4t9XlQh9UnNX39hmldFMISKvVrYfPZ4wqnMatPIcxssl2agfOMB1hEwyGMwgkblr837XUhQf8i
5IGvSrIIEvvMNVqgEIq3vkg1DoU2DWFC3l2+Ym0rEIOjtnCDb1hwD75zynJsiowlbesDP+QA3Gkc
UZr03+H56V/2ABtleAPHGrhm9fSTASA8ItYgk5HhlAGmXrMHItCAqeYPT322s3kx0G1TSF4EJ6xe
+/pKjtfsD6Ymt/gQ4xLKRCSe10y84A7uiQD4kRT2JbiLGsjOTXXbHjzX0fn6w7k+qDK0aSA076Jh
f10YxWZYkIBjOndKgQJRRWK8Qq5m2e+7cnM5zsgOTjc27k/MqgVu+Son/NYqXzbeODqh/fWS7Xsq
Gi0sS8v+tslgd60dJaT+z5DDJPwvyX0JCmKPtRp9w3CWdldeybmW5ye3zrsFw3VFDoiHir7NNhTX
PIqRa6Nd9Xq4QSv4+d8Z8qKI9DJzminkM5uNhqmAPUw4IBeMiP3cGaytttmxsfuTz5RyFeeg2mim
kSwJDs0wgU3A11zdFBTQ7bUC9pl9T3vYUzfSQRVi9YkIqzuCIMMWsPi2fAuSrI/m6DK4t2eHOgX2
MCp/K8mWxKweh4c2mu6MlGJt+UjEKzGKriv7ZiFoGR9h3NmDVJ44C644B+lGQKO7I+UI7ZCRFvyb
Nsyw6ALQWErcwhStBHf8AKw13QmC87Fl3KsNQ9nJuGc7ZW6an/gNRRLjfj4pzzOz37usyQDhcz9F
KMyT638xFoqzHctdSXz2iTVUKdP+si3xiP/KHDcV+7Z2VILJsXRKiTby2SNe4dF3og1bsfFtxVjq
rlUazxBPaXQfYnq85c72TfQEHvhmgFOds73YkvbYpgDLx99caOhLCqBqbhU8hmBJuIih4jEkaSBO
gMbAYlbf5t9ZL2cy/ZaIrWB9EeWWEkZ/mhGSATE0/+lZoaKWoMI0hVgFkkEdyqMHFyJGpUaxq0R4
invFQ5Q3+Y8Ll9I59WYe8Mv9i4Gl+p+FDTQnXbtPpAyeybClGS55zNB5V5a8WAPVvAyXCcWwdQOI
nc7FLvVZMK22CnMlUcERW6N5maA0VTGVoqFmkEgZPCXOelMPxuNo/uvg1gjqcHF/3ZTOfTWi76wJ
G8naj6+iH3z7eCBlFbUwKWWdo8rfyoMi/oopM5OHyAaFzcfLmObjrfN7is6SB0MiDGDmXK+Mf0em
HwKAT0kX5WePik+4SBvRypV8+JBgMLyxG3QLX9hbFPQS4whyxURqYH/AtiVcPNTg6tnf5UQ9/V22
XspS9X5l09qb2e3MR0EC4w9+x+M9iwyquOAXu4C67v7QfEcMV4+wICHHYIwmGUhh7GZsaZJ70liu
ISrAPMVeLcdyvArc3MwTI74YZQiw9vtOVqFuF+LX1W6vyiehCtVLET1ev8pdeVEja6yLfn10T7cB
NgJlsNjaYUEB1CaHQXb432QfmvXMDUqdhHxiN+5D8u9nmVq+wxbfcjmKzbBUHkIrVoK8JYvOcQ16
+CwIe8b9ujRdoy82AZd9eKqFudiY/t2NNeaGPuL2kuJejMDIdO8W/0dvli6FAJ6SPdDwIP/2HQfc
nie0YA3za44As8SJmooI6tt9HkDYNcpyi5sDGFHVtX5/e8sRWY7uXN+m0tLV+tOZbCUmj8P2pqZr
QQUXJ3y/STtLkDBHuwWVfDc285myTNOFll9Z1PWOYTe7Jk4D3WvbCnvusb6EHX6Eff6Oqq4r16Nv
capnnWP0+zjzK4yaU3bOYpRsPdA5fylj07J3iig491/78S9VGlCajt8BKdw88UXlx3YfazzeE3Ww
aoHm81IqflMhnQcXXDhMI77y1QI+1Y9Xl82dBayHPBWJbPcFO2vauBbV7lEwi8+7Im005PTxFIOm
REeeEQ/drR2Rk1Eq+BaHNkmVKRtCTac2aip6AucWHBOCjtNWaX9H/oQNzaMRfux2IP6QbLIAjgCX
0klz+rwGZ+N7TtR9/FfGU9U2/q20CQxiWkntOpVYJKC2b+PXGqeRVKeeFv61P9EsuEp+c072bnYg
Id8+KETZFtMNas4SW31G0ifs5uzycvvD9zI4mduLxm0mTYYX+9jTeCUccq1Q3Hx5LDgMClXmT7To
g+E3kh0O4sZeJ30iIX1jT+U0VrPOxOlmn6+3YGR49oCbSjhyg6Ajfq0ojGTQ4T5UuPiRECzIV38V
dOjBrypdVHKds++fhYurvF30ixNWp1fZCLs22+MDzZoz7jH5CvGae0jJlek763TjPHiZU2/VVauO
N0t/Fx60dZCbTXMZjf1HUaioH1kWDsKXgyCO/Av8SEwvY36TwdQZYsDnp7Fm7e/zealzrVL5bwel
ocwcJpq9ho6qOh6lG6Haq6RnRzDlcciV/qTqa/ApIYiALthKKvqkecJwzGJNvXPUoL3OKznA1lBP
o6ltZ79AHXtuPZqX+orwO1nTmz5QpzOBImyB6+lt11+Etof5aSytl3NpLJGYzcV6tpaCGT2E6zcS
ge5Ws1DxKvzgOhjDMA45akdnGbt6XQL2XpuOUzobhWKsHBiiIw7IF6thMeNWPOAEJHNYL2pggvug
CriXRJWTQNoDEzip37QM6DIzXhReNOgq+NLvAx2jZ8caeRRGih7GN1TNtvaaKMCIFLPphnrRD1Pz
W6AGSuRBEYPqxiza3XGipHgyb4ZfY/s5Xm/Pu2Gnkzg/1OAst0w6zikzBvGvwFoU0Mpw9fjtfHzo
M5Dh+cwxSZyR2COnkTv02wdQ5dvLNNg4BZEg3LeOSAjl1IfNWMcca7HGkbKJ2/MdAHLH3lSYyKDU
e0QHPluPz4DdRZ8CLQftv8TgwgHHTYxrtrwsoSMtNNRyoXPRrCsgU3AxAU1kHXMhjC/fpl8uKW0M
BgmMhYFU2ypH1Lun7B5BbxcSO14rE+N4fj2fmQjt46iXuo+pHCFOkFeFYdsVk+Ss+TJhPlf0MYSi
k8sf3IqkIbXeiiYcvqVMcyepCG+l7tne1N7AgJU7FYLx0y2VZ0DQLnv9ZNkSlJR4Mi99P/1qCUYN
j9CABMMZ+2yc1CxfL4QjE5d1t81wE07LURynmeJ4pegI+IQTt/m9RmBU8+qUQGmQwaxWsL2CtR7d
q2VPYz8xLjN/tPTnQGux9pWKegRsEHIz0AZr+ArirVncXtwS1YVD7Ezdn+wFF8W0MMb4tWRFzc+l
8zxb5Fy3ywP/ViNZT8toTsFRDu4eCE5rWAWhdDsgO08qH/KmWSxJP5XiVA9nXvp+KsBHFziYgkHz
grex5Ym8aG7m/EjO+gJVxnCTEzWZrLUL1p6V9NWOlZbRFjCTtu72Yhx6abE7jNqveNHZsbDdwDRb
XBoaBJ7kErt0160+SQczLSjQ253oZGOvBaFQrL/y0Gs9FyfrR/PJb/g7/B6SdeSdKOzHQbFpODMu
scIXk4USHqXmY50MWhDE9XOJoUcjAHHhAUpYqoG/MhGtf0lhzTaaMD91bSs46WvrPYREDU5mfT93
LQeXcrtEtQ8hkGHNNUD7jKOkcBhA0ehEjc9/BVm05+6iGHe/YAlMXntBEKWgpb5KcazaT3y4kt5L
Bh8gZN7NxsguD7uWJybulIJQCSWMy3GY27FM/RKPf9sJmtaMWhqRRzouKqvTN9q9w32YrMW5NJZC
7595Fw2u3YFl2GP0Oep0SGnzvzNRLVImSdbI5jZAWPM0fP3sRjke47ocJgccGDT+KVOhibH7PVV7
CcWMJox4OoZS6cwBvj8CN2KJUNcecfu+9tTfzm189yWO21vRoBsRR4oTexGvn/cPAtm7xGTwkxvo
kSKAuH08+onjwVq8LdrEorV6aqhe0MqGbWYLWu3WKiIA2o8Xim6bnPmX1p4vYKIYnBtrbMVXzQ0E
kL9vEJwvBk2J0+JRFTpxAhxt2sZfzKKAPLxl1pmtGtf0lbA7YgF7NZRLs0Iz/7WiqqujoQTU50B8
/2YrhiwAFSK1gdXEdqqGX94hZf0r6NkTngvsjq90/oRsVQg4/f/CwGTxqT9roa9AlHG61hHCISuP
K2BDaUpGohcYJMQxsa5D8LoTtyPN8F+Lj17Q5ob5hthT0PrHuvZQOnehzLl0MxPYprR03BvPORJ1
w475DSBFRsqHYhDlA2h7kvbJs26lo9LuBgc7ELRcflOxtgSJHASi7+tuVz0R6yrDJma/73wGG9bo
higScOk0N9NnIdMiAXx95mzHWOBz1y7tHMUoK8l7xAwlWeyq8DegY/EbVcJmfBzCAxkwTRZpvivv
cihmFw71CSHyu9Vx9s06XMonzSIVO69jqNrTYa/rE2C84ZY0Ildx+wonfiTvH2aJ4KHjxeczXLC7
1GVptUlb4uH9jRrbuRVQNpHWOPfiaQxkU5I1Eq60uGGBnGjqo3wR0CRJi0zO/Sh8XYDCaxw/z5K9
SS6OuPuRr5Q4wsWEtsh6iPvsmvRTk6Oeufzhr9VwkSynd6BPVd5JiTSHfQSjK3q3u+R/Qu7dUBXY
pbVOB/nl408bPIQsf0TbxknydRfl26c8fvN82DpD3rbn8gGoPFsSODsHSzwDOgzq+n4toj56N1jD
2T9+JP0LczBCjJP3zI7yBsnl5EVIw5kI8PIEX6lN4oDXPAYbB1RJdMuLfcbqIoW3elsWikxjk+q0
k3US/ZhYuWvekOZFcAUuohu2St8kbOndzjoTml9//+pZippjObz9ZI/kT7p0BhUb9sufkdvADz/U
s6R7HNNcK8FKg1tw+eR6unkyBFK9WFlxPooqd1Gxvlws4OZFI/6RxqAvizkK895WTCV/KiCseeH7
mvxb0NKdqeq/WPQrZsUdbpaLDR2WXeKR9jGRadi5kZc9sRQFd4Fj2VqpN+auWGy5rRSEm/67ievy
AG+nIYdPsL743sH03UDV1S6+T9TFRP2GYaKF/QtWWvVu/yBLfQo2T8aR02HhLWWxbyCn7wjBiagP
vFaY+Z3T1dV8qVtLpJ5f9FY40vGD4WmC//PfF5Nu5N64E9KktDV6XNS9fEQx9h4bQ0kf2+B6yswk
nchQ4sVs7VaR17xRAbtzDzQDiy8ygFiFAYcsmi45vZCLyyhMgNrrLg7ia89HDmh2bhFmRNk8Q0ub
JIwYVoBO5ak9JH/uU4Qt2ZzA5kcSzvohdvz13BjpzXKrihhsQ9bn4S+XGUqNKM/FOFz4H0XtwI9o
fcm1GLAI3zk9TuAl9DRb1mJvhmbdEhWq8gJX2/MIl1eeOh+yvLrCzzNc4oktbYwk6rW950C2R7L4
/YHFE8Pix++p7BWP+1FN7n0Y6FjMOcMLeCGCTNPlwyfb6RHBNGrfNMpQHE5iCQvGDdclm+leZP7S
6CZIJJeDt73b4H2Chib6M3LDWFw+9JCbR8XLqtTu1SHGMh3+cKxqeci+S08ShPJJxzUuz6mlj17D
A8yuSmPcM5/e0BkcrDtc8oPyrfdBqLhd7BKjSl5TEtObFIms9Y/V5fmpVqtK5EPbvYV0NmLPr8fL
MtxqLyMYqZhc54LSo+Upj5iJbl2dYO9tIYUcPj62QcQZnhU0KUJjFhB7gmIl2poCaAP7FYszXjuE
qnV8YN8pdo3Jc3NPmD0p3gOHrBWgbLNhyzxWlIiUwgpjuwjDY6AnmWkFy5friMdh06qF4UjJdfa8
huqgkghokx/ywWSWicaYAqBjFo7g6eWS2X+M+w/6fFlPwlmOL7N939t0ywn+975aw7H2ssZZt7Wo
gZZB0tgrWhEUDf7yuV3m8TbOoRrvdkefhE+v/l06hkuAJqu+zcqH+TiqXgdrIJlFe7LHAoh+doxZ
rBCLDqETVabNEaeX3zRVrmXm44RCp4wtVaQbSLudxnlYEAsA6WkGBrvgdBLRlIItmGzWhsh7bQae
F6PEBcTRG+nIBTYvuceOFQFQJsO2DK4mBXgms7y8OwGbGix0gn1yQWoh6TnqOTdbjAxQPRqwkluy
CCml4+oGbdBZPCQjpmHP2XjOWW+PEgldQCybeTw/w8vv2cheOdOTLFt9gpatmlbYG6T4AlNsmouu
cUhGv4WfDIivy/Wpi0P3YnD/vqa5M79W/lFPdY3vPVYsBaQQfLmx8f7KwAdb+BsdGpvjOgA4bM7Y
uKfs3K3tGluB1Kj5c743Me8RF/GaDB9giSJitsltA+PILYkEhEwtpjFMOZ2bQf5gxOXUTJ5pfiGG
u8bxJf0tNo4mQ9uR+S1Rcv5IadstuSpaMBAl10eOPVYC06iKKsoo5zlbzB69eiZv8U+LF0hfGzBD
EmFwQmHz861PO1jZXSSJEY7vvsMUC8rKleNExHnyts91drYNWct5RwI7i42OtEcVPmC+DkII3+2R
cSoiI0ruWrMZv1mhZQ8UvEJ9FrKrOMBKvXchGeVBODtg1V+8hXwoJCo+kEYvwkLPfJ8v+4Y0S1E7
9eisQ3HibA6JJ5g/ZKoduJwVM6DRa5Prks+azHp0gj4ioZuMxWjAHGxRNN+O/vcjHqM+mhtrLfJl
4YbAXc1m4Uq3435jZCZso26P2AZqU3/qCg9LkRtQnrOYU92JxAgJo0rmi8tC9Koo/m73Kf6VjaCY
welllNcqe09pG8KW42yzxdO9LhyNJJSKen5r0Lxo/BLO1LJOqMObCEbb7R9joC95FwqI9JhBF3zv
9MYL7r+P3nF3ycbEvoDpf6IhbD0oNzj8eZ+tU51RD7jp2yA1yj9inaDrQEptEv5tsms4jPqjz0qQ
SZxnihKpexZ6Rmb8w60bXRWK3nC8BC3SeUfJ5QeumQk5sQahL8mX+ceAmFSEw3XYuDzK3SYqz2a0
EEpTxHaIG6TixQDww49CML5GpFmi7m2lNzxCJZO7yKVuUnMnqSTSYXsgscjTZzGdVnEqv/haA0l5
92wlrP1jAz8nTZh8kkNkFxleiyswbZ2Xvni9qrblf4LA4zaIwTCHo8t9YdxuNI0uSoufC6QR4MnQ
Gyi40EdZsjAhyrvk04DCaPvwv9K3vrKaPJg2t4suCU/iLVH7webHcYh0qOZ+DoluAUD3f6vp/FFw
KvsoybCJ1Sp1YlvyGNPmAMU7Fdp5hIPZPHVL9kQP2V2DlEMG5KocLhuc8yHvbKNpNveUMI7ofZ1S
DN3OthB8R+7gBoWp6/jBWkw8Jm/WsvpLMrsvAXhPel2qY9hdaF2y183PGMYiyiUu8fqNQnOX8d8S
Cfn3qVI2DAhvlpt3oVwy6gMLx39b8NXCCU19ADcbjYGdsacj+lFIrpfna0HL9Jue5CZOyee5MRnD
vGppVvfT7T9cMz3n9Dcnw97oy+psUcm/rbZsjEh6AvGOxYGIAUyH/3pxeWz97+yU8pC1RGpGlwO4
PrnHc6IqoFYvYzOz8rQLJuUWCeuNV7iKkaptzs2eK/A6B8I3N0ZgbtIgHVHXK0JmTok+IvFk3lGP
jTMrXfbrPwo3oGQvmmzLJgBOCsR2m62FJsadl+KMpq2X+75AJjrqRP4wq6Ngea3RA2mA1KH3W3YG
ME9ySP/E0qaPkP/d3SfA7UV1pv/uF5OtxjmViSA4kfQhgIzaSHPJn2gY/Qkrtxs59ZFBX3cSQ+zK
GYx3MI61MH/mMoiK3A70w63iQfTimGHPpndAsNQNU9tTMONCdCVvWUDbX0g/T+a8/LvS/jJ5MEoX
UPzCB3HlQmP/Lhoh14evBkQ01uKizd9Z8GqfnrJPPtygPPp6oclfu4pe0pcXh5iwvymvf3CR15ot
4ohEcwDLtIpEpXunPS1WAPoD4Hab3yWMykXdCGOwhcSNN09G7ia7RS9VgtIIUDQZbNbtxNvmEC+5
eFPhrUSUjFmlb0+pO7mlLijI8vvZIqhjFlQRy2AELwzLqkp/Ju+iJt0hYO+ZjFdWMcUBSlGHT146
rKoi/A1RGlhkJNGi7UTM03TIB5bt+mmvNuiYHzKJNAfGJoj/wM80gcLPnw1Z0qzmIKZpttI3nqa4
dDdwdL0Gj0+Z57dOU9n7np1Oz0tYTQBGKzNfYK2RN7sj9Any84Qy2cvL41JOxp1jvgrtM1BzkcPQ
m5OwuQ85K5XvTt4O0VCmsOkUvcQPOmHpVEAHECsGzAR9VHVoMyB13r95uIGpatdTXgzfKYiQlnvm
6O/5Zx2KxmxGGwBN3NXYOTRtHb4SzyIeEA3k+FqpJusV/k8Fl+xCL3bErR/oVUVlx98Rkg86xeI8
Sl7ZMQ11app1zkPFkvWL0VKlAnzvlJH3X08P3sqV8Du+QQ8sWQ7BgajiTClbfLMDG2KSZ5WVU0OK
RUyGryWCoGMLr7tYrIdWIJQZnYi0KRMebCX+Gr1ANyXf4EUVVgATVnVYf4KT+YK0dVoK1PQlksTN
g7GnWM/qIpXrrLsrU0Xncxqhpp0u63lI7Z9doL7Nhs/chV5zE0mnVDhk6g+VWRQLsJfzjJ/xX0q+
WINzvflBY5xT+lfXdWFaSa5bXtfeLe6HC9ptp+CKgC4Fa80r7w6pJpIwJRrUCOYXn7dAFbC/yVBA
5t1+Ilg4zFaAKQY1ifD1KWg937gMDMp1eaPO7O7JtDhXynvRzwC/gMKRJh9CrfkXokV/axT9PPaO
pwkc/PXLyISoLhqn7MN4i5fmhm2YitHGD6uMvnxzXINmezCGnTD38bC7Use1Y3qnY9DrycePsG84
YN8jM6QaeNR8RYVXmv0PeL3wqxWpL7rVV6LHZiNp/Ye/kQTg+8X+MDP5gIiLppjT+0hldSwLg1Y7
XLz359wBhb0wS6JyzK492nCSdyj3TFzRBpK8oxbSr+TRCFfQUoFHjwJPQreHl8+iK5vpCE7DuQwM
MQ5rEz1e3J6FEMR3khahScZlplRvArX4CaY/Ew2kWyHs0ljZEPrresciuqMVVtDDiWeFWpkAq6h2
gWRu76Bo7k9lpS/WG3WfKSI3i/XILpRo8oeSeYzdXG7kS7ezMXR4oGIDwjB7pfFElLrL3RSgwW17
P5VqYU4KwwzOjM6XncNeOYTLi58cCy+m8tzJ4orMclzxMPfoeUO5QG1xZX+D/1pJFrMH56q7CSdK
3FNJiOEllyEQ/eN90Y9hOLPthqU/GdL0VGamGHu54QoDu0CBAc3mwxADfRaIAvmH8Pz/FrqUW53E
dIw1jzqPQzLvK/cswYc0RoqyHkLLl/wUSSJdFZZH3IEIcOKzFGDdugBfxMBB4ZrQ1UGzHtH1KG2q
hvCITdMv7he9dOdUqGA2vSt1DRnlQPXRESNz1wJ+Ty76Sv4XsIEtTz2OBsanRFB6jbZgnE3I+rqg
cZn/jHgKYfJO6P2iTyLWA8xvPwESurVo8APjlE8nizlZw9ktEa4pAC2F+dt0I6NBNPZaPStqBI16
6dgP3yBB3xTWMBgW+G2W3U+t7OaPNfZE0TZYB+cGzYlXSJn2fdMDp/7ko3lHcoLIGneNLRO/Ew93
i5/wFFyd+IGUDlmdvSYQOXqGNC2XsPnYTE3JNIgTg1wqhSjRFhlKtYedutpoyivXycSkDcZxaPJQ
WftuxZtiG0wmBaHT56tGVMdGkLjmInfQvECkeDJEBhKJ+dSzy7dqno3JeKJ096IeoRWlGjZFbqcw
qfZYCtcwEJUTVv703I3DAXBqaHREcld9zn6JoWBI3fXddr+OwpUqvceYyXeek1Gu743D4oulp/es
UaLWXJbl6GP3ODiM+yjNdxdCz+O/wscOjcFwU0cBuAn5a55eV25BTfxpTEOBqEZtGwWESxzTDKTt
ybKvOSaN9DHwC7kv6ZRd01NyCr+XzU/znfy2y8i/4KLy1wOHTz4NZ8zF4s6MSmehzwHcOnPH45cs
NHkaZhsz4TNnpncrmvynKZWthFesSzsqIJmqUkSpe58omPq9YSagCEx3f66bSuruHYcNRjj6Xm1T
c0JeyjYNJ1ID5DtyUf8Y41QH1ryj7xE2SDFLjvmtZEsGX8TJDQ9QzkAzTTLWh/wHLRHw/53Y7tyS
0U3RxVCp+FDJkTWur8DBJzzVdo43k7W9YKg4HOG6zd1pCsmjLUwWkk5097lhKfKh08XAlBSy6mwY
6wB58iX8AFlA87FpUjzaaeh7F2JKdjESl8HKQUppOZUtzxwM3NeajYUXsMOGugJUmfxxLSRx2Aas
+VHoH35FB6gAFR3ZAW7M8dHXnSuY555RsVLq4k+SAYNQXdtlZp1ybpacItf0cWQAT9s4XCDs0rv1
rTUPeX8EAKZBpy6hy5/B+u3lUYwZTPmtaEuaW6PxA0D4dHAKbPT7S8ZnN8L7kzXx0UcuDqYNPPU2
H+jpMmmLt7jLuQdRYhnE9RCkTIfMvlb3jPZD2nzFlNgUqbxRyZw+DEwCQ9sR+gbBnoDn2ZYWORFx
up6jTTJd6ruP/y6LfjoObmNSuC7kU0gyRNxZQBv4evor5SQfPNvzcKciyuGCaShTeyCCxJiA+F/G
wgNkydWgNNI8taOmy5WTuTVddqZDSUXEq5gKfC0FWVxBd0TYQBRWVW2nOU3ub3ap9iORB4ZFaaoC
QFWCvvVo60ehiKNDydV7dpDiJCVWqZi2gWC+Fgaz4Tufh8SOphIwijpEpTZbMB8rp1n3zAB+aSCF
7C33Q5okgOqmBzK1GASqTm5aCDOEeOLZtrlI4cUDaRDRFq2CFw/WAo0mGDa1TUgUEGLsIxLF8/QN
EU+z1xG+SHJeA4cHMgpu220jw5j2sR64k+S/3cMkLBrDY0PZZmy3v0iJrpJQ65vnzmgaDyJ4gvzj
tAOydsYMdnFnJpy0iGocoMz1m92MN0yYvp7eK7pjrUKg7kRbm0QhbfoVpYO9n/+ySTAsNZX2H7Tf
2NaOAH56LesI9pB1zqoNDMiSkL7edyZvD1GEbbYd5S1a6CTw8IQi70iWRw6+JIyAuDlAnhy3Zyhs
IuyVme07d2YJIgFyNURtawOxES0uKubSyn3ZVTbAKaW+596gKgKpFPxeRbH499TrAz+9LzKwMxz8
oC/33aBM/HikzuZlxQFzBJEzaTiuwK7VfqccYd0NKHnBbl52vBVAsgQDM2fy+Lo++Z0MO12MqX8c
iMNwDa/TsHi6Eh8pUcbB0d4G9GSXQTsmnRpXMxhH8ezUljLbMuaOdBK/paXlHwVpA2SgOM8BizsJ
ra+yD3psg6FGaMbyKzAMEABVFXaa2qqiQpXtipIoJzzEbOmhNoSCUqavKEw1GIycBrXAMd7m0eji
xVVTyaZ1TJDzALxNt749mv1j+SoH95Uv96IZ/XZY0V+KlmcgSfwTVS4wifBp8RCUrpKX+eaL/qA4
YDPUAVdxFBKx0DGkhkZPvEmS7siCq4opEzsHVfZ8rK7DKUchLgHGsCtNsVvbsEroW67k6SWCQHB4
rdTqzQEBZ+0UJ6Vt2ZykAEKH5IiuHqsNr8/y+STh3tVdNCryg7USf8C/s6JJSNF3fZenMu/hwl+L
H4RWMBpEZHBqNdQdSSATOqq7W0ejnAYZoYTeukEnmQ9bibPnVMJPJm2JvBHN12gF01eTUWPYbHHM
uhsBwc/8lIYtVOoQMsAr86S2p8uScwpyzUBxOMKjmXfYdXhXNrTkF7Z1MTr4PYXeFHhc07XoXJx9
+F6Y6QAxpvF5GHozUY5z/OQDAXDpKDlJukcL0UzyUS/lr+3Gq8yRLR5tpcXWn0epw0bKdIrQPLNq
+HxQsfyMAOGlzGOMuCn4IVNeB0676yuMK0rfpcYT9aL/A3EeggwAHAOb2ET+n3AH7TLl1tHiZjIF
0GMBwjnmkrsYgl7gQu5DI4MHWe9PxUMpiqwhk/AOWmdh/PSSPOq0gu5nD2vCZTCBqAB6lXr2xXTf
XzP5bpgtV2scYdCC/TfvF0axiekM9RNlUNwEGTDenOjVH+8M8HHxlDP7zYkT5zYg6qAhz/14EEFd
ssZaxMIHRUYRw0eaD3sZfWn4QtwPsk/z50HVZDtJch7f6Y/m2ZPlqEeEdplYx5Iam2eo0qlVmYrP
IBvwW50e+EH9FGEUVm5dfOBL0X99/DJeDDXhT8je/btWyzO0m8DU8znGxtlfzurnDg+145gb4M8e
+vBacWEN0XTG62NU6cNlH4i0zfjnavaTLSbdcQjWaoizub1dd1CGYGt1et8TPDXV/Nruzm9S1TK6
RlpVCkRNNvxOTBjJ9nizOi5/JhLkZ4IJQ4kDGMhgoggOXwAxw+YnOcc8gzEJ6OYi+k208IXt7x3V
pLZEztNmNcswIkg1sx26dLPJNbpBAO3HvQ7kvHVE+myjtfVXkpf7evUqrSd+w38HYFmmeVVRV3D2
xmvFvTp+rtZkKREY7xa/ZmNAFNlOaL3qSCH2i0y7Mg9D4CQHO5ooPoL323bQ8yBtAXi0uOCiT+Xa
GbURrSzZAYtvGubEA0QIxjDDDSQ29VLnbcE40p/uPLjVW7f3r47VlW3tc7uDJJPnJfR6FpcodAvh
t15HOPoQQp45YKUxKd6rTvSIc/rHz90Jnu3P2/ieqZi6Qro/3pUhTi61X+5oVGYK6dF2RaRSOiz3
hhKTSEvkvwaoYiyZYsuFAcS4a4k5wgdldyECPvzmhBys5fmTBOUMFCWOotlSlTqhRTgpl15jZXh1
4CNuNqMBD/aLFblpmKyzNcoEbDX6iDZxxiTCSjhfGLF4w+EEntQEJlFyworgPKKOP7TlpK1PQuYN
Ezmbc0ow+U5ZjofmtaGfG6GMei30nNTTQUhs2kfFR6HbE0aAFcgoxskOjxQoP2hM+aBNjKyd9DBb
zgTrYmOwu7ZP/8n+zNUMB/hEEgml7dd1zNC0LIP3pdcDX4pT0Mc3iYtE5fZJ4hCZNK19roAC4p06
YjWNxuGYmYXxyA+vXHMugbs7S7yOJEjwymAMbUnewJHJyUg0jbp2MYasKvmMS0mqdh/bmUCAd/UA
hpDHsyM832aRTb47VasgfV9EPKEOyok3CheCAgJOKHDwcDEtpdPsI7kb9VC68ezyTgfQfgMMuvF2
1o6wpQBAkVHJZZa2dhtwEIZxn7yzMf+dRokcoyYY+id70+8wByD0RfqC0Ene1B/P3NcaC8d1tihr
9DclUCUe7l87mUXVU0lrAp8ghHZe3DXXWAMWeuUf6BiXFgyZx7hdUjc4M/XaJ2z7X0sTQ3VBioKV
e9RUGkF+xVo0vCAPaMg2YWL3hfhhi+qxcn+z32Hh6wGOm++3ctkmZXxc753TWnXxYiMc2JZxc/9V
ugM/ZwqYTFwReV3v6SOtSIr+X5fDvt0lKfzISmU9rZ9/yr+noydGL9v56D0Ie99IjQQmNSUJuO/h
roGkAXgfv7NvmtvgrWau0aYhCR1/56l3TDpz7Bg2PbRz1MD6a5adt5X01cp9aNZaoZV+rnuQtUQD
mio263pi/29Pe6M0GI76Smvs5c9nxhwj4lrdYn+xgJZ/d/qfuyltKdvgpAUzBCNKMpSD35HW5dTX
5V2QK8DkPf5g7osu4jmiCIdzozzNt5AkoRo6EcVl/vlSEz1lqiRDy9xPw98ssfXuMaQpYODBKleF
0MfhGdEdUYYWviQ/OTxF0yVqZoWG47qozvk+aFNOup9Cia6AfucRDPXLe68jrVIPQx3yqhGbxh31
8pbhIBVzHpdddCfQnvLbrZJ6v6nRuo7IeL8yWcsTE5GMMReIzgRiM9p5oW8qvIwRCrpwu7tcMspB
FX40ibgi+awrVLgi2YEDa8nj7OubvnszEeFA0utFTpgmuMBwJSIoBnvaR/Q/U3hj9d1xbFELSvLY
ECUGXW11HSY+8FgsDvdIxHNcOEno3UK5x5VzxAK9um53QE2/3fCVFhHqp4sflaUXRFeEqEgxnNe8
slC8J+Bp82Zd49wqEMzCYj+oWE6Kf0P58DG16zd9oQZkKHKUCvQMh1c358vV0qe1f0CckbJUqRIv
vJl+1xtaTTGKyT/xBsJlW9TjJI0xF8gDOvANe/UL2ZTNALMbpTPwYMdGR42rg+pY5OrhUlIRzZ21
SaFZdjIGY1wO0/HakoWaAvu08IUX6miyfDw+3xjusDCWMlaBkWM6aFhvHo9GJOIC6etuKZadCv6c
UmbCuaV8y9beDcJsV8Wi5p1FVQo0PX6l4NALt6bSKr18AK9ZqK8eOJ7Mw773vXP/gvSX5TAvvMSN
sEQnTbypj4l7k8oMfM3sCH4MUt7VNBU0Id+LYBN/poR9CyrGP4bv4S3ACTk/LwbBHfrVkvRnvSQh
GyGAe87mcfwcZM29gRpxgY+gViLVasmbKtt36av69SP1Ta6hCrylLtOFmI3pNrVGZzvQUHfDMy8f
5vgtDyteu4Xp0/5pqYr/NNmitBnUA/WnDQvTXZhA7cVd58E9p32ScvJ0FWmetojRjkQGXnN+eGsO
dIFHVRmt5xCtV+7TJFkLInDutODC9z1Yu40Sjh+aT9CN1hWwHVwwaDFV4cJVX90xo8C84/IM9FRJ
BnkAMRv9vLGSxi1Vlrb26cEKdk1RYtIl3Jb9o0JL23RdoNfmjAuyvLgLGABrLK3eJs7yZNM/7cfj
3FC7oUng4dsGKBfFXa7EoZjhTsLVVDA60ho1PwFyZTC3ZhKdS4SUTcttJHp2B6QChXzhUtcobJzO
rOZUpefbFbf7qcPUpP5S3Wzv+r7oU7qTTl4DooMefoAEYU9aFhfl2MeOFXvXHu+Y0CC7fXHtkpgG
4kJFotSSzYqlrOjb/7PtnEPV9tiI3hARtr3CxnQS5c94S4gB+NQqaS4vaXMoqjUBOf8vyIOO2HTR
MnnlrWIHhNTT31ScQsCqgoyljCm0zooZoJWihQqk3cQWkcfELwbulYA5IfO0KrEdQErPd78h/XFr
Nj4FNx0kvIxdYQMpPOsU0lxfnPLMo9Mnn1UFH+I5X10kV2XGFCbz+PexXbR+lxVsj4JfCgnlqN21
waoLIQz012JxZiaPpIX7fNtQxtO8PGsSBrOd8RVRemFKv+Tb/g0ZppENELqVXCTI1duTd0ezzpEx
6WWxoODWHHGu8lK098U3x4bloCgeMbSH9LEpQ//roKIq84cdPMWtqfhyb4sNbR8RzqmBlqXLRayF
Cg/gP2KUJ+jHLcnDk+/I6Ypa6y8t1A2UEXTZkWKUhZoJS2NoI3RBJGi48kh1U4R9zvF1adOzw1dd
5ljJ45x38jjMsutlndToOk8EGVX/5aOgJJ6nyr+g/y7MYT7kK3bhvZfRngKRm11HczYRn/Tm565P
E+jOQjxw8vKvZE6m6UeP/n7bIGQ2yiK6lOVscJv2Ezh8QGkpGFwbcK0/at0k/3qzvCCByrRelYA9
UpdJkzFt6NH2EwK/1hxDya+DJv4sjVuY2Nb93loTKgHpyb+fWq0pVveXAzjG0DnLgO+Ppi3sB9jE
xaySYp8APy6aEUPj/wQ56kpKXnRT82VNbExi+PkqsNGRfoZO9Ka+tmZincCNRWqj+uCKO1e0/79Y
erD1fiJ5vn5Thb2xBgi4Fbj0bUh5olRA2yA2DWQ178v0kspyqfzDUS2usIthYI1MFwSmYFhX/1jt
qLiRhbr+3mlC5PbQbwy+6p0jJfTQF7SIcW2gOuwutXAJ7rC6MsLRvmCNfsd3wJh4JlB3lMXqUp3X
9CHc9Kpqls9tXqKb3p7CoAzSqm4Hs9X/atZ7yRSKfJbYu1dXXe/g1kxuwiB+HV6AC09ClQf7pgMq
5v5c21ov4Ij/QUnw5PEAJeWlXFwtWIR9mVPeGLTczObdWtwgmCftQEACupuX3oktReNPR94RE32E
szq8CpaqRaDSAQ9+WwtkGsXAp/sg801EBj8QA/UXTFuLGPQxJjoe1pijJdGEneaYEUi98Daejcw0
pCA9HipzhEYPjsePT6mAV2D/mS1Q5ZC4cr2SFR+7bZTWdgSwSY0ZNrGA1WSuo+UAx7hHsvXr8gcS
7Otz6a0TiMPgVXbw8arnplVR80lUMrmgmB/FupK7WRSsl0X3i2X7O60E22siJKNrkn60uG6L3Y/8
g2AUri5a+HBtgG9uWp5Bn8qOkHwM+q9nWIYJwknF6RqyAiVG0Ca4yR7AfviQY8Zoxa4AfL/HoZNH
qW8LScOLzWeho8fEtg3ZtGiV9o0Cc03pog2HCbwKQj2R9NG1+Vs8pts0CSWVwMPxcTBSXWTD+mJd
JxYyYpKMKy3sHPRZRfYII0OGJaqqctwQjJ6EUlqaj6UIyJLbIfMmjUoEvTCHOoHKGBiKBQBvXKew
pupfdQNbtB/rARjvX3E4h+K97VOfkno2gqzUk7ziXgFngRO0DgF6mrXD80WmMjirXZvVoaDW5nVI
IR6905jhnOPNZqPONwpfDDqP9KTxkl6Hxy35zW4qFLk+5IW7+Uu297ww2ggcBgLXEbZaGbh7q0t/
iNlbisQtGd2dxmYtlhMyxSaWlUsQl5wy9cW2u/SLND44jIhS0p1rUySSuI7qqbQI6QibWfbSdhJN
AgrD18k9zP2fyabYPOIVloh6yh2VDJN+SapDUcEdxAcYtqIMIqW+B9RczKruBmJJ7kAtF/myvJZ8
3kgPQchEl2GkKHq/MwTDchhS0QThnIB++oL0V9KbpIsIEqbkqf5OMXVudEJ3U7pvr5AnB8QrwN+4
lS7qYiPFWUemj3GLlpA+jrwOO/sVbfNwZSGv3U6xE/NyivqrW4yZ4qiOExLes3ITulJKOwuV+Gfl
YfgT2c/jiiioPI5P31csxdk1L5BuijRy/+mMHDagnk5CTJSQRSpkJPg62l4bY+x2g3/rXpgxJzaI
RLeLCaegDCyVdQR/TN2MdaZLZ4A7s4zs//rqId5DS09lfqFqrEqSzU6IO22AQWF20kUbOv+bHGcr
po7+W4MstHFDqZpukfJZEsXbtH0lZ8biJTPKpzB27eay0MwkONTLOzsYS1HyH8t9AfZxnf3GCbkx
ymA2j7yuJyyUt9tlZlk+0B+lcSGd0weGgcN2Db6NCHSS4aR6EqUw7ImM3acSUmZyc/rJvdcGR+01
QevLvwX2f7WVudXldzJTy2pKn7oLl6ycEe1cUZYHcE15XqnbAPPF2qQuqFryOuYlyAQZ+dHnCaOh
g0IHhwkIL8QyZOtOwU0OBJPz3y9HlV4A1olESc+muj/n8O7MP2ucG3MUuC0ijOZpXNOzxIt00Z4V
LK6J9c5qhNi8n9Fsc1zk499v2fsPdHeNldfk0OzTwpdp276krQxItNvRhM5dpqrZICyUA4e9igNy
rlDjY7KrCATZwR2FH1i0pW2GpBx8wKy74aPwYxj7lyT+56A1Ar8SdUqjuQYfhdwzpyBpEAIN3Fee
g2RTgXw2KkeMOKT5HMc8E5wNLU9JUuJvzNLMs4z1XOgmlFCwlRygLXpEEfIish2xGnFi35TAmXeQ
O7GKkeiK89ZVITyewkj/YnpFCIYXu56f0bPtsldXe9n9Q0L4nxIs+kMPdhBjqhA/DfZ/9V8V9GSm
HgEiXeFdzRavvijyZlb6UzGtz6texGVQYjFFQPxNv7irkZjR7MVBQOJmJ2exuRu2cMN47ugizIEv
ofUB+Wup03KRzxU5uQnAlFX2W2P49wZk/LlmCCwy1sgVbMj0Wlz4dL+FuPuoIASioLiZDEnv44NC
GjzvGo5gHKfFcS6xZ5WVng8ZI2FxIREh4+D9K7tNMeBahdma2rBgh4PnU3HaKXhHQiQFztWKAiSE
00MW2kHgQeY7AKHpm2M5n8+fAvJQzhBOCurQXc7H0d8NtmUVidVFjzj1WJA+RPyGFqiRkNWWLR2J
vg3eIpSTdBbDEi6jC9586yJ+bP8+98hhEzyThFzy/znKkfVxiDR3GNTZOmHvOEab7aoCSZeuiw6G
dmuo4/HfMUmXsblCCdnCZmHyr+/2voqtNsbKInUUOQKdDVA+MfLwMoYt9reL8Z61opoow3qAd6yt
FsshhJHvSRkDF4xu2QV+xWzOXMmY8VPc8rLNI7faXrOVLAWDnJU69aP70BZ5hiREXNImvFzVSJxE
dmNdOjSbxeXJ28LkWhuPa40XLFDkUiPx3inKRRNgfndLDpSuMIFfVtcSLCSLFOZfN1JrHqJPAoQ0
pwa0D1411lV/BZEw+qjQiircIA4uKm7AnMwu8G/xBKN6K3u22WcE8DhrkGLNPAQGlfFg+XTJuQHj
C37/fZMnmbA0usAjoyVrZuZLRyvykNfzqDLdw0Kjse1PIzhaGKNXdeaK4dE/ZyC/oDK4PqG1xZJ+
cB4V54DPwghcl2QoyP5CgAlA52tNMb19NXYMPpUPzgLqdwOI4OZnBciH8afh1mcFk6+RUgMphvef
lPe0dtpR4Bv0rv/1cL0wIniVtRtlDI85XNmKzERYiRDESPcTG1cu9j4JIOn7qCLIOHGbhD5k0dpg
LauqKrI5vVHN09nbmsppW0buDQ473ixpDjXoIfcLj9lGcq3FL7S3B63b52YbVq10inInuYYvReLH
Sjz2Dh3HAuGqczi3lpoqn2w7I2C8VJd8HuZ1QlU7PHJsCxJcmuxjTxESuTo0ck64WMvQ6T30odFr
FcKjZpSMJ2wFPMttX7y4r9gAK+CNd6cFuvDpeZIWQlqWVs7ySaBAkuWCC8QZwNbQGGi3ufonCRP3
+Ug24GJSp/PPPxk19CZq6e/x/6eduSC4RAYtCSYIR6sZ9c4SJbBpp5UZkkzhmSFBiCRed9qLkLXN
SnEcYLT0AkMuKZva8Lc6gGIov6OuIEhUKi3iyIqnwae6ebgoRzuf4NTwu6qiFn2wVsM9ScYgHsre
QnCu3IA4jwG2tM3OUaEnGoispwfq9b9KpMfnUgRFpKakliCBQpru8AQKmOCGTOdAAQDeSimbsNpa
qI+xeFJD/OWEJHlzjJm1jaXwlTtUUTcogrXeJJgqeRYmMo0PQGtt8zV5JHyJshANMJESyYG4JWfh
K+Zi6PcG2df/Yf70ohAccPmxSBJNjnGRASiQDCIelr/TiSFD+awiNHyV51xdvposIb+zE6cYak+M
dsm24myIrMu1Blas9QVeFMWHURDdkknhZxyXxG5Q3AlbOdvSGETa2VN8CC6EoEvJ+WB6LFDGS2zU
eQyLImlYge+d1fJ1AxbVvqiCf5R1SrnG/CAPN+dIYFx9UiyT9I+bG6SIXPCgXaXVbthDHEaD94Wy
nUcKX45Irq+FwS09HM2gW/lhOXNbOV0P1of0lK6ibNoJOBd6VNX8JrJjM2LClVSv2njST+jQNveK
+8Sf4RcZwFsBFZnLY9zxKyek9+WOONEreV6UzXl9TyABpl8D62QzZUe3S+Nn5xup7N8XG3dXR0O3
y1w0K9N/tLDr/XXi0n0vAJYfuhRO+Wemiip4u+r/2q5WqokkPnX1y3fumbR+JPp4ZLwEZRRh/mY9
U8wDVHTyE3yonSJLIlwF/qahF+DAbRnmOiyWGeLnf89kSz1IvBGBwVqHMVuIXS5FMOhR5CRo1Ifb
r+THRL6YywHIm/KKUrMAT7B1qu1zunZIIpqVM2c0MU/jpctAE3hara+MNOPSfrm9mQ71kMVtIr4J
SKob7Od3FgWvEDWxJujhYVCcC9LKtroaV2+UHa8mUNP/CSnLQWoTeaKI+TKxeuzxjPETvWLILGbv
iC9quDU/R/7Y2mbu2V7w/X6H0VdQKujov6JsPVesv3IYom4gGfks70KBjA2cu4MSH2o+grIJJRVk
TxOp8ES6tWnmEUzQg8pKPUuWVGOCK8AUWO3XUarOmxOp9yh3vnE+Mz3GuZTUOfl84/nEFNQxaKa8
Jx5/cKtniijZpfXvhus58d/esrE5bjvbWOyRdRxjnWe+e0ebxq9OBGlqAkB0uAfXQYASso1Bh5ys
sjI//dBSItURq9J6UIrUy0uF/QNyUBPAPtUH5PM1xAZIUjMoYfhANvVnccUQKhjCDe1x+RK7VGor
A3xC+OMUJXn5w0ek6wRn102Wxte+f5uFq1eP03ebi/IdqNTvCxPt92UZXqn/tsLl56mzbX3IZfcL
3ElUKbZqqQ55qHHdMseagEVkYeu1ST4Sbj5WTrLwrcaxg8IbbpdzimStzfiOmIdjJXuSHpTvgslr
JnfD5s8Ib3UWx2FrQqhGmVCLq9S/csk8OCzu2Bd/cnxwl/SjCumln3V/sHkixsRz+n3hknuZvrlk
vXhw1CwBqHFF9LsJxo7haMRGmpLz+tQyAkc+CM6VP3xaj9yr75ozVxsVPkAHkMrkz2TFmIiO3n1Z
caubQdtjapA4sQqGmxGMTiAfW7IYuPdNCJSeNRu7sKIBpzQ/8Ga97tn+LxRBMryTDSujOeErKCE9
y0qhltC5X9Wg5FNMpZRRW17vduwEcHhS+E/W6q+tOyGNByLbhVhit/lOpMHZd4eDNWt67a91ftWJ
FBORD/+Di5un4UA1ximFqVs5L/Cvv8jkAI8mL8rCDgcELj/8Qcs2E2DfulXUoLgN/M9xl3hLfaTi
hbXX6cGswjZAdEDJg/aMaYHHbMvhO8u2oKNzKep1jDLxpPLdwe4KvphoqzK3rMvK2QgQ1COipLbo
kgYsNdUoYW9sOszlfoWcLHwDzqwAwhsv1fcvDV4DKGWo4nKNoAT0rGtlLgcbO67ZbttAFXiJEG0I
cHVEqBZVdrOUblkQ+kgSDe6/BmXhGk8Tp9HJMl1JmMDAZi0itrJFrf5M14zL0qp1YpqYTynvYEB1
pQI5sIS2tL/iiNNlmnjSFaCu6fFNqSUA19qq4PjkfsTYGXRTgxpul1w9BagNurvyYf/QN6JFIfVB
R2B8KM9NXMsmspr1IIwawtrloX7Q0FK4cErNFgcC5b0JUOTA8nH6e++MQYCDF4MwvQBMvFlR5S5h
Ga6H+5KgJrRncy7WAkwMWMYILB9fEYr4I/pjBKYGSN/QdoE54dm2YgcmmMStx/PMAOEsg74tj6Ce
CUdHHD1NKyQMPvF5j8uqU7SJDmeYmZKadYBOUVipAeMKDJESTDlV1TUKrc2hml16nkjK/+BUxnGA
PSHtflHjUC7DsxstZPlR0SnbKepBtZ75qGcY2C7BUjlf1KCa1yVT/VDfRoAqHbYeKl/ELCyFhB1j
sNGzUrlzEBWYgpJ7MjxVCdXReKP/fCg1xffOX/dfdEFXJtNUiy2CaX5pDm3nZ+lOJ+v1jafTphH1
12qn5u99dKqGH1Jz1kTL+zjWA+/rQqwVzc592nTOTElfwxciX426MdBMHC8ghc9uFJlHyd7gyaJk
ac1bSFtWRS0fzZWuyCzkvy8ie3XojhKzaHXB8Txf/LiZ6yagA6zDLci3z6tnvvKfMelj+laMXt+i
KgdBTJ0kEH6zU2Yun4LUOd+KZe3zdh5fFLIewy5Hbblo8yKCvjQ2oZewjwCKG2LDzOTcDa5hdmPn
deOcjAnCe8V1eVHMFH2ouCRQJgKGaxlCuP8+WqmiusxNzVwiR/7kRvFRnb+282HHNjz7ttXFnmZ0
84B0209xUD2vLavQ60Z028rX46DMn53vGjZjAuNj3LBPgUzMZXs3asBMpiduUvCrphyUcb6yxjkZ
p2O86NQAi2czGjmc3Yo7Po7npHJC52JpACIgJrF1ueMIAEZMqmUADlD0YiAftvt36Pv4M76HHjxO
39sTeBpmoHFvDS79QpObPx1ldggpwp3V90lRkQelOScoV0BSdc79ZiVBGS7f8km9D0ySMPOv690H
MOxOt7Ok4bJD1zKyeW+VeAGxYQ/BXhncNm/4JJINNzfaIRRmpHL7LJyOKMZxC75sj36BqTSjP3Ur
mjMwXebmuq39exGU/0P/2mqiNBfKmaAgmQAhExHM6azrFQILSGuT4s63wTw9smtkz8lRtSOjP2hh
j+vMjrO/0JoButpe4fUjqUGzsEqi2jGdNkPxwwQ3zxoLodirbNghejyWD1ncvmb+oTbYB03u0g62
uXiXgAetRf9P6wecTltX9mzJv8+W2PYLf/VK/WtGxZUkv8weOni2fEediaRrg+COwU545F21wBTl
Sv11GwpeDRe+Cv4Tc572rcN8ZQ+gV6TdDrXJyxcK7IAG5sF7Tm1fU6Zrj1rtG7nTb6y4Yxf/uXf7
mSsDczIzwqUvxRSbFffFMjiDCi41JHclqAqmTBJhEO3Mf6u3gw8sG8voboHmvckBXg+ZJKxkWw8G
LquI2ZZLoOMAvh9YcjxsuIDgsn6Opeyk81aWYfu6WzI7Gqb/yZDwup9xWbnGarW1bUBnvTRga9GT
HAvQXuzFO7mdRomJF+jtZyTRwCm7AGX6fzWUd0oPx/R4euC3WVhQg4g/q+J3eor/KnryR+ZEXH5Y
WS9FOxwJrWH1Fc+FtLqIf592hcTZDzZsPFKMGHqkDjJPyAUdcbrraAfWlBUU71oYZCsQ0ptU0cj1
MHeeHumSUqomQQPgq/u2wdfZ/jxAYmNh/9EkuwF4YAtVVEJZVOCebs6E7QQIUHXvbfAROSLLuTXq
k/X/lSDYh7JfNz45iOAcfz2W3p/D10mDctBzbKsyJLXOSO/NKhv1USyIzshCaA48AIcAJncNqQul
sLK/q5obyNYIg28Pm1HVEF2gCIABJUepgbO9/MwdPHbwRw1zH5eQ84CZeYNyupFtK3dquhaza752
0x1JWrqASrutNUSBHYZY4q8dNCdY0AHjy4aLNmdHgVAUpF/yipg3W9CKHLw5YAFuQ8U18V8UMkq9
Ox53viu5pgRan2faif4HIw2oIq6qD6KPqEoe0Iu/WLDBd2muGIZ7a42i5mY12LdXNa89QuVQXUbz
nfoaalyZcE2SosliOUjxGiJrCIxGxqSDZtACMchbPF8/2qn56OOcmHNHyteRFbm/QGoaBhxtwCUd
JZEwq9t55J31vpYCBoYVAY1Fm+yxypC+kwt5ru1kIyE5SxOxGGTLc25u3hOQZvuFbCSc0sJ4DmbJ
08DOQ5cy4n2zKKEXKTZ8ZKHhaw85yEgLvP5XEMkCf3I1Ea3smycvSogslzpCeJy8U0lUmcuXDFu3
UMyXRrGAiuF2rTEYY1IlRncIk7o90kuIV3KSTqkDCiGJUUZQ7Jc8XBtFgsud0R8NCOgZ1+Xjazch
n0lnUkTrkORaJTrzkhUp2xlcR2Ak4Ntp63CNqkTF4d1ykDSY0p1Bm423r9UyuWN4iqgsJ9tsoso9
pBEuieNjFmfTm8LgyVuPDXe+pZU5d2EE+MkSnnLMGOSJAFWda9/QXVqpMLMJqVf+j3mQD7uBZSNV
1uCBgACJPCoURWJaeSSVg9VmnMrU8xB44kbYNDzA5RqTNRm1kKetTrykSmPh1TO/N8n/oJc9TpXq
cn3+NB/QkXZZnp/Us+oEEXWcVBmYWg2FXK/EzxtZMoey0//9mv5qONzMpd2XYNRe7VFQ4pAvFeNL
X/H3r4/w61noyiL2yTELw9WJTPavyxRRvoh2g2Ia9uCaCOa+FXrwsimpLFNxalQqLdDchXsFqvrW
VPbIZMgYqAVA4+3g2iMGTy0jbC1oG/JusIsoDaSLiEGi3IXrNKlu3o0G6bdKPpiv7YqU2IIBl8lj
7igl6ZJFDFyVc3vh+UzhYa8r/23ptdDissofSzofL424T4WA387FU1+RsEqA1D6RG63cSrEf9+64
h1/KaHr1dP97B48G1WHlpES0Ci3DYC+CyBxkWzouuymEpi9Rim19ZVTxtSUmTRrMzGrx/qj5w0Bx
KhpwA6gBvab59msJB/07s5CEb7Cj/DQ+k+OPWB7DM76cMpNG/G5Yr2kiUE/8+/dFhHeqYUmVVvFj
rPZO5Hvc9quWPGyklfvIJGM8Uz/5PzoLXuY4EVqlerBCT6mxi04Bspf3JvBBTKtalgeiiRdY6vO5
V+k3ey773ffXKoYHJfu1he8U/GhlZAY63v9pJQx+r2pNs8VGKN1z4VtkxE/Ni/KRZB9dbTvgKJ8x
X5kqNmttYS+ENDHdKD9FfymG4RJP4SJTJhiICY97BjRrC1eDiICpLHUJ+rzZsHhCWJLrlQOlDga+
hC+vWU6jsa/1U73H6eYxSWAaxotxq6hJxsl5Lv0+7oA0RkxDzHflZIBfu04s+4kcRkIn3Ln8iZtV
/gyEGP0lO2QlybL1lH3yIrtfI3So4NUq88iZawjuWGCVaeEq1IOfUygZLc/Bw/J2sDDTJ0XSAGiR
oGVCR6f2EXFa2NgPxszFMfIEbpH3XKenapY+wS5g/TCaoMyIplch2eD6pb+abLM9EvtSBLpLhS7T
5XMstzklMqUNckaJmSJ26i18lIFTMlSWZ/k77Sl173UB7xsNMEf9U1XsGNPSkyn9D/OqNqQbXotC
BbIlgLlR3Fc08Y9cbWNnRDfi9rgABxI7HoH9cmQ58S3uPEVHl/olE2ERP6jNAlKqqCpzdEwf/Uo3
pN0pkmc59Fx8KkOsULuhzfXV5dxe4fIa2hh7wyX6rAN76LpLuSP/3LI6tELZ+JNSbnQ/5tTrzTOE
xRd/bsDb48UfNOZbPVHo8U9912Ht/JQY/naqzkCDiqrFrzDp9KrqO8Eh9eTZhVmIKDeoztXC67aT
hdaRDBhu3YQanmDNU64PkifkDyP9mVZPQbRUpmIoK0ZpO+mVgBCv+X4S7AEzqFr1Xv0hHiZAheSQ
LBhEVpBLtVx53VaqtrxMDLSnDLICBVoj1ZoFYxUk4HVwKs1reLJMP++DplKxd7YWJoZ6tocIXII1
iy9G6I974++ZINeZEQRU5qnGW+toElXyMObzyaZND5y66O2cXMQz8di/oJCBzjxSwBnQsb5DO56W
CFSmKVxPigs4A5wOCpJGYCGLrXHKMcHdPBSJ70yfi/BWsCOpy6l7VpWKRuY/k9yWl3W5yMefD22z
zymq7HOgr+sEdhmVbIQunULjiwniNSrWnGrQvUKF9ZcQNch5nmFe4Qi3/WhlL493qlDCCK3oY+fi
V+bgpUdFRJnBjEkHDJ1l/qQBTTsMevmi5arSusfn5DvBj8leSrygazT3Y2pHCvinElKOc1vQsRle
2XJH1DZMdVHPrKvvpxD11cSAqoFfu1sLiZwFEXnAdRqKnMxNs7Rmiaqi8+BgDv5pPu7yfG+gY6P4
YuXtApJmv20G60wgAVNxlH817pacij+iNa2QW/a8hWS2uhaYXQDgHrz54WQ/BifOS3YJ6DcRcmQw
vshXWwF6fAl+gdTKJ0QJCIyXBGyuP6AytBKMrUHjdHZORe1aWC4izG0PHhFHVpdhX8FZLlVZ0YOO
EcY92Z2BXBMnJ4XpwvUd7Vxw8v05xT1hx4/1QHg6JqxPipCNq9XMJ6+dhfVLt9osFgME/KHt9Vey
tdSe+laMny+YbIS6twdvY4Mz3D3PxIMTYRVrBtvOBrKc9KgR7/kdB+UsA2KjbLqCj/ewwiMOGjkW
ofoDjLafxYCI6eu3rWwOXNGLhMCmf2LU0+erMyDAgBUi1KnWHbItA8o4+wWtJoJZuENC7ffeEUlX
luxQ/YtTzk496Dmqj1+YkczUdElhZsy2m3MYVogBoWXtR2mJ1SnFCSp42OXoMnOXfm32aurzA74H
RogOqCs9mTz9sY2YQSlGQGrpBmGCII26pyje8xmjQgTe+IIPCoCFyZAQmoKK5b1JXf4IB5TQnsgB
ZsCpvUhhDpwX0Ji8EJ5dK3AdlGAhUyLyQlDdYncBvPfgs5AQwO//h2MOByZmlRUn6l+UN2HXwbkd
wmjEGbuuQ9kZruU2Sb+jOaaUInS/0cFTWTucosHryxyvHGFI/af4ZsA6vwDDl2q6gCpuqf7MANL1
hLEQhKYlPupQS9IG0beiUYejahzjJ1nYpRgVAc192HdDMf8GhRY7TLmOzWoKfoLQCFevm9ukizHo
Y+0wyEFd1V1NfguRLAlVvlAtF4jMf1zbLie7QKdQ3eJXRiFc7sBYNFRzqBB7m7fTFgC/Oc7kPS6y
TvWuzRr5NAD2h+CAoK9NZ7R97VzxM2HJxpW4ixUa8/q35M7NRRXYxwL2qO2bgwXhFw/EbqUJZJLG
a5v8jBosmJMvslB0oKLnFulzYgIB3osYyBxw4DUNBpxcCXdj/Xv/bhvQ/EKrhw9bRQkV3lz1ZMf0
AvPJsUfMmnhcT2uRw1QSkw/Nz3hl6M5gIk4DaxIFXoDgMG5Xkh+oqfk/nsCMDJGlSBktvpjDIN5n
R7A4cAq2dcT3CDG1NY16D0zMdA0zs4gyrI2SU9pEmMpla3lQX7717o8a7Lt1vlf0scjUquR82iyg
P83ImyXAJAd+Nn7F6/gj++aGnAPe7H9vP2+0oL0eYKyH6YIFi/BcUSlAD08qUKJoOmHhl9D2bbTq
x8cL5eoPrAPekcqmZGsKLaY6AjrzmdS4vAT3uPtI6LWClbl3ypqWCeskJD2+vK3sYijr5jGGiBlk
zRyPKPb3UpOfhF2i233VZb6gD0ss7IrGkZiGq1+f2H+1fxl6qHBaTUZMuovIaDOEXGE8wLUhwWgX
tfheiYDjVXO0F6L/nzxU8B1zIfzxpXumCA/BLCjzWRHx9aSMA16qjWl2ASCGksHPUck5D90NIbD1
EI3dsexFr083dz7gzfcDMPaVUugmL6Ke3Zi7t3FimdQsLCmaIJRzGbEJVAb/YY7GjmuO27Fjoogu
WGxKlzBLzFWIQjVuxb04/7eYumCXAUK2lhgMJ3WtZxiJ95BCJSSrliztrT0+2waFgXZ7W5+N/GH6
9PH++HrYLZSiaUy+hogeQz9TLcYWpapRuE+v7XqUC99odsXox8R24tfamjff+p8/97UFrGy9cNVM
XZhTPW42AG4gnTSEYirIFt1G21CVLls5SgKa38w/Y1dQlnqAMWcOnOfVXFs7WcoluxfAgqr3epSu
68PMIOlI1CCa/EcyWJs/s/ftgztZWB1U+Bd4IX8QMthaVfq3ramh/26aT2MNsDEJCHqU69PGkgY8
SFpYR61FeEVcexj4yhmaJhOLLpGVeWL3jn16+bEmOiqY0B4vNy1GOvpyg745uDBNnmg6iNJ1RS32
FbeVRgyogHreyP1MvpyPBFAmVHGXZnw6Xs5m+2VhLMcBhDH/KvDgJ9NmbuWsuhGcVs1oLljqZ9tu
Ktx8ymPBf3y5OSyy2H/X8vxveDdHXkz8zeh7cvWSkrYEpuK+xFgQRilMjMMdEwPKGE0SJXg7brrh
x1aeatopPJEcV8l89Tdw3dBQUqAei30yhMp4vQ4Vb9yIcSoBbuolxSoea8hPy+4ylKcWnv1ANlOk
QAQOHvIrWLms3tGG8kB+zu8h0/rEdu81Mq3NHXhr6G+LZJIATsjAScM4gEKKR8PZ81c0/V+xHEtY
lFFEg6vb6n+/l1qLOQOK5dfs316hGkTAuT+ktIES50pd4Cvcxp1p6mMXGemeyZnGF3aCF55OtcrY
m90aI3nHAAv8VGxFt7pxNLk27jporW3FfICrTmiqbGKofhVgugABWybXW+ZnAGYt6ZcunnduJ1JM
RWRWHQlM+Mv1tmFDH7S6AvKwxY+dg3P5sASzv/R9nGkJ1zhROPXMd5svNEQGcLWNScJGVJpbygWj
qM2xI4FZmBFePzzGqQIpESMkn/5cwo8QtvoywzaYGJxoBIFW6MTsh0kPTlQCzJSirdUbibIXJECu
8Y34cjg0CkJCzj+hTREI7vsjdFogzmnmm2oasr0VyBKNyLqj/3izX9yBdVo9+XSpMsGHwE0LHgEa
MiwQVGQtcfHqfNllmr0uQ3duuP0JabU2VFU7vQOUQ9GYr5TlnotHy8tUN15LBaIBwTrTABlMsqSx
xeyWGXQN8mNfHN9AQsQJDVL9qYjuwyl2Hy2VEZn4MGWjjkUtjpE/jf5eeKN0s5Kd1P9Glgk6VOBu
ZDO16pUGYbEx2M1UnOZyaNya0VVXA95ovko9ghXNdx+bvb4X+0XUlgH5yu/OcReSXTQdjdJw8B0M
vhxaiWPgaG/D5KuR+fhQh1Snuyd18HPcHDelKx7aBsHIgy3Jr2gFn6YwKWM763UI5dqOmSZhqbOP
ndSipBM6xFG/0fqN4mDA3Zqc/KFz2eqwgHqLDSEWC9D+t2Tit/sjdVGbwD9EZGygWGeVvbOFMih8
xAiO7I1GVlyOEGhglQp2XLTb4MId2xMXt2v2RD6sMOGtHoicb8LnhCWYWgWubbinBSiXBQlCpJFo
WjuAb+S9Gh27NilVo1b3uSE7uVPUmiEIpKKoAmBCkT0PCIiAO0cdlJfQ+3PnKlHa8egFrV44hKeW
hIb2SRZhLA70LmOMjJc2iyQrNhgLqCXwG4VBE8VP0w4pA6WVtZjq7x4HnrQvgCNS3LHIeooOX2aX
WdX/PhC8MtDSAVov5SP+8cHEF0eU9aTb3E0/mRuBcb6Uweu851njDKCqnCA62Z35mB+MUqutsDMW
EHKQHDNWPhQbqRNDwsrNC1F7BFcdD7xRqqYWfIMRe6dibOkp6L810q40v44Nxa/LiN39f6mfonOf
r11M6nsKCJd4otLN13nRbhQuYJHKOHa6Yvd4VMHK4cbiEukeKvoQb89oRZXaERVXeilxrNtjgWxG
AnvNPZB8zBJBFDNl2psYA3aKi3YJILLW7kB7rsLS979Q2Bt3StEDZqaAajEl7n2sUofFnv9ejKpR
wgz1i15oVJQZvHhCg5naJNlc8hDKD5NJWbaYhWXKlFUu1J4UJFoDJ/Baj76kVWedEKm14dI6hB1x
MRKKMMu9e4J7Sc+JSl7PyFGrthtoVsZxBM/78ixbCTpD20uzJ80fPNlgBJAXexAqXmNmrPWEH5Qi
J8yASaW/5t37E96cf56Y5yq8qX25DveMegR3T4JQLy+ZCf1pASBRV23ig0TacCdHRFTcaa6tpxNA
JV3IUhT+4kR3cbttFmF6EFJoE3BSkg2ehgW90mcqDRM8SxWaX2VEJwnqqmzqAADQxJjupweseOn0
76uTmt8/MeghwRl8wA+SxNa4bY/xmoCr6P6FJbV4bdrUO508xr4TIoQ6EO2JmJAjo2yOWWRYwRKe
o7NGQJlgtWm0d6WNToR9biOn/rM5aLurPXjpoH/WIldbvqx/3g/uQk7BDzHHPY5TQZNJMpp7CHhO
2uf9rznqHIA6acFgxVISfXJhPOn923RJ4sWc2FjNd2Xd2SQNjZJKxD55pnsSyffpxjbWNptN+CER
anBgoZ+cP97djge047WsD08SAHXjvbww5EqdwrwxuzFusPChITil/tLW/xxulKuGcPb8oJY1n4kL
rDY1XHBSV1Z/uOwyBFe0rUpXYKaNskjKQhDJgwBH+yGPkxzTZRVQ7teZaBBc/0JhT/MTxr0SPYzU
G9AlKyVbp2/XaaR945hj3hKx1DGdA60GAU/kTXlJ1GnJ+AHEhHEAr6qSM1tGgNRjc32dKu1oPI9R
aCoXBGrRIK33XyOXscGyioINHqbfzUXKvVZ/2DqwuVEe4Xd8+XdeIeu2ubeBTDkNzgvyEBXYKH3P
6yf55sb/z0ko8YCCuSBqZzxHmaLE/6vQNuLQbcvgixzBTtTxFjMW6cM0AXoh8wzzJhjzgCtBi2We
8myJosYxedXWiv4gqJ6+dUq8hFRgjGWW2qNNOkGTaZVGE6zldzPqOZ4D1BBOyZJVEeEZtnX1uR7D
e6btoKIOA2P6ZAikzK5M0UYI+PxhhkVNGHjkL2zUAQ31eyvRXc6m4e0ANqthrrq8Q/xmZLf6j4U/
GBotoBctIvMDLE5+RbND+8hG+ceroJ8ocAMgeGEhAkNwWPlxDKmv/rXwW+bREqnRG6PWnFdDiRkI
bRWnR3zIgDN6OITwBbBmTm4s5QyFPakHwvOkTfatalxBdhbTWEOFlUPEmINh1oZgB//NiqNxJB4v
4ZPMsvgCDe4TSV75yLp1UNHh59dB/K0HjVApVY5ScxRbSeekbqFK+cji/ZcPyGELJkM85PGKjjTw
IGjEby6XKYg7KDBVT0X6F5LCHJ9FsH5uffFVUGkeTcdc7cHo0Xcg80bwXbFH3rRbRew9lUdmh4H+
Eh75lp4jeNNSBnH2/SgncPekj36oqZPxy2IYPjW+xCJ0H3ur+/tCBGp1SygT5vN80n6X7iYIRJol
A2t6SXE2QVRR5EVY9H5NMbUY23zf+9x2sPae7z3YU0hK/RBVRbstUmtzIGTtbSqnnrSQoTH+Wuz3
wBKxfnbfX90DphE0PrIvkxNfQqOcI6VizTpfeppXxpex4dd/WTQpkF1SFFBb/n/Sq6eS7qIvpOQT
vQv8foh/IN2segAECPLa9UPs/Y6+Y5oSMS5VVUfLo0i8BaYx9mfskxkdtwWtQJL5A/YW6vTSXsnW
WgBmyOiXba9Q0wM3ecnmhSnmeMKDfQhgK4AZTupmdFwu4nlq7C9A7Dg1rgYBXWVcotwMr7i226wq
/Ia/StO7qmeG+ZgsFOvgSK+vxqg84pbVwNeGrGieupc4OVi5yipuXq4nvKN0BzDjtSuOrG04i5h9
B6lT4WXtV2afgOU8BAjPj3Bx/Mfa+XR5SPPco8dTq7tktgt+YWkL7wmFUjU0yqDOiAjfMdKJxoAO
XxTlg69UkuLD9A4B6cjbcFXP8/QYwqAhh9MZmuKkVedeZVlStKF8fRX3eDrA4Tdk3taXDG6TNZj6
7Iju2nGm1lD75MX6AxyPe3JNYmUuyLR1EoY7JNE0nHHyC4zMm+mUw4/za7RHJ0r4gHnunL+J1XQv
xU11E9s7UnSawmtmBYWoj3C3c4BsJ7ZJe2tUg3KxGpC5vN8Ns2rKAjdMunvUxuKJiRIYdjObeZYH
kyN3ymYT8c46S4MkpD795bh2nDO/dfxbVfWNTEHgVtksvLPwhGwD48/bvZ/pNlNRxoArN/il1uaG
u0PC0oAvZOqZimQT60YBJiMeKcnmp5N7lVoJTNupW+xVpcty6llOUOLKeTLCSNx3+hiubXNHm0vT
i/fcHauvlEwtuqq95Yc9WHxodkUqFh6q9ROOd/rrKfcsiWfyrl4q+OFvKVnRNXPR15tvLsoL4xpR
ijQlANXFOkSPkhzdpF5O1a0JihXmjigVm1413RHl9sPAX4s+oyeDG45lSZDIYCPpA8t2pN1Sas5S
bMEn73yJRXwP5CE3ItygNYEP8Lu4DgYP7LNpAIdgnIiJBo4u2oEptNX08MiUkkT+smRwyO8I3YBG
x6uXBM7v6rxYYasHfAZYqcUzVQcWyHq/arIh23hQiVWAVLFliWzBKsbjgAifocA8FC54MLGOEOav
oIbeocGgIKZbmbBzQlJo12Fq3XrO5GPV7J0hY/YC42Q8RXEf6DKEOkWOwp8WRY3rk/kEJHlTpl2V
NWnx289uYILvNo2hJI0uNCzBEhsE0XKP2BuJ4e4HwkCk7aaHCm6572dlYGjLuwxqEj90tpCHITc0
gr7eFQ1dbvSRYj6YQjwVdrgivlKlN10xTfeg5ex9svKASzqhsWGioNN/6DTlSgswoklW7tA+bPWz
CI/Xo0WCEQFQodfpYyI/faOJv4m1kTjaPZwvd+fxekVx36pdoeRpEErTnemrf4C9JHd+u9a/Za4I
zIBcJuoLsCpXpskAIErX4BEueb0Y5wghcFdrv3yD4C0gH2Y29Ny8A1EzR2w6KusBC3n9bhxNq59m
UlOQLNY24nGWckN9T5bYgYB92BwrSbzIpmncOETWlt8AMChGuIJU80uAIwcz2oc0ATAnwdHfEEhZ
8b85T3XH7yyPIojuHKYHBtp1MHnQ7LCB4GQU9F/4o4+rK4lg0QLBK5iWLWub/ajRDEwm5yXViWxn
LW1pQE7h/yVJk2Uq/ZDpe5jtHFHW5BfuhB6JeH/tA7d44TSxAOb4+bkrYK3SpG3j8zCUQ6Mg4dXv
lDgLRvtautGCHJ6xHf+HI2R2qoHUeJyTS6GC4PbFEVhKyywQhshNnrmWlAehWrcLnMaiElMPdzMQ
c6FWSBFzDVvdcxNIvrhs57HESmd0z87v6TbYC/zVFjiCBohm/bcBcn5B+Ls7pIlz5D9i2gaKxUOP
yXkHQ2Dr8Slsn0ETlSEFOH51+akkIW2WSeC1Y94DmsF5xO4UhG6e9NTI1vXBuCzuBOkP72nE5+vq
JIbFO2IQUeTHk0DCAsCFfTRLqmueLYXeM67+9PzGi18IQSr8Mkn8b5t+qECYjAV1I6DbDftrFUKL
IwwhEBTcMqLcb7n2kzPzldn1T72qqGtHHAAFG/ZVHGF8CXl0/gpjtHTMp4VKCNOV1f5T8oqoiar9
N39xCeLy41cQju7a4sQbYDeactYZAo4pxlM79h5bGATnpf8GzFPmi3cwkfPhjYEeDbhqW6T3Vv9R
E4gH6+2QhFvGTzyk4Z37ETp2ByatKKLbabpq1mgwkMJXQwnlkvH9a3H/N/UdvxgesBLq7/ExWpfI
yjlNBQFaVkXPGmWKx0fgzWyzAkOzoqeYcEI84BCDtZgi9ALKMVaEOJQqAaL4RdODkGNYLg05AVzb
lHKS6Y1wgdL3W0/nc9Ks3pX3sWBo1iEwEuhYPkTJqsmZbiTBVSpSdAIsmBomquvSUXy+aeHzVAgB
7VFBGGWJVDD8et4jyTDPjmIzOLyCU6ql8b/IcuEQAEoKiIK7ZFsw/kT5ZYQQDYVrWpShAo0DFh9W
0oY2cIShUBg06S0mZUUWBAYVp3SeXpK7HeIZeHkT5E20aSlkLdMMJ4189WLsGT4u6XPslpmhHLfp
/CNwoZvBh5/eIS7gsOygTn+dCueaDI8cTKA5pj25trE837c6UQgWkCQdZmxDdHdO9jC6spudyoNU
GCvI1IC+ovGOFVQpXphBWnaOFS36UoOENTHK6vH61pG6zaqBtwJjlJyNhay9Z7rY/AsgQrmmgSvV
YgCLsEsyccwAqUd2SFpYeL5wuPIQORmMZ4D3j2WV6f2xxrxHlyA41kYfEYogUmstUBGOeg46Ho+U
uarAtP/ru5HU9aN6A9K1p6UAIqwIqhKJ9QUgRcIdBIRqULO+HDOWbCZZ5G0PeG+FI/NiiqCLGzWy
supwLFoFGCDxiIxIkkmyPT2oe1CVVEo295+10BcSN7Eu/o2wpl3qp4CIQ9RsQMQmmK/V07ZqGWF7
ZDIfoUVS1RZVCK68UcFxMLs6OWHY6yaRw3TxCnHGAJTm9LelG8xf5/qYKh1hPOU3W1Wl/Ip6PSEg
/TM+trpL+jxwVrOnYDa8+BXRd6aGYj4/IWnMDkIMWC5oVfYwBEHfNNbfD/hquknRl+2Vf+XVsIQc
7SEn2Z/xSfP4FBs31F50MmGP3U8IivlyGA6WTs3y3/EUtTAruq3enq075CuDJr1eoEFBcTANVo+d
Exg8sXXFeG9y0FDOFvs1nMQWvg8LAITNbqSRmHPidbkYeNsojw1Jz4l1V/49u7hGN4rqrlfe2Whm
AK7ScS/FwLVuE4JyMdyeCkvv+YfB3zr+2PAC7qNJ7D22B9iZn5tL8aSoAGBFQTHl7h1b41DAn0eu
MGkJqYMhBZb1AnHFcHQsuoca879/0hmTuOGW+U3KFxEzl6LQlannhyXstP7Qi5uiA+JWDagcoC58
PQo1MuIjdCjKdCeyU0+o89MAcah0A7okGI7n35IZ+U+BYweLjhAf0WNFW4m0JocsygPPAEocRZIJ
9XQ9XklM5bjTBEPHUbYcoHPzkwOtLITPDH7k3jTHJSYAXvN2T/0z/2qCN+WhzSfEfkZgXW04E1El
1xgyyvdZg2pbNmK47iUazWeDfdTU4dlM+HVNSq2MkyvDzXnips53HIS13PzPHiNVA7mbwWAQ19kt
TaSgkSU7ew0KAKjOAp2+rs7c3Lzj76ashs75YSxkIa9KLnhCjL6zX1lM9u5PelWFfKIjTZYF6+xf
GtHNByqZZ1bEgrlG7baKWXjyXgOefAik8zg3luK46qX5I2+XGq6uCEluUdyJ7/+Koj6iK9ubDHIT
OE7HJTyjWP99WOX0Bm/P/vtj9bYlSL9e64wPB5qsnBQgHuIAak/mI+p7v2cUTWEczv2UUSvSn100
Ir7IEfGOWe8c3UzOMbeNIbhadBMzNIKnZbY/bCveXsPz5LLJrar9WFm0Vov0+IFsXcepHyGfh+IL
rra195rFgaSVf9bUgCOyxFrfntmGiMUUn9zFoXXzaxvGmauHrJ7RNHLNZlva1I4IMWysY+tBAHrJ
GzcA/rKaKmOCux1N/J3xTca2UAtRKemGUqqYONsDcACLhD/XRDVtWfDvXKAhv27Dtmq2ogTU+T/S
Vvth4oLf5RX6ZPC0i640E2dWYQdlrbb6YyDTNbo8JUIiZp6MZrLTBcGP9Sjl8993p5sflg36xtC4
LIFo3TxAdIjvB8DpSwBSs9OrpwoGifMTkrfI+tLGTqT5kQkQJw1HGQMqbKPVpVv8Fw598tHnIxfk
i12tQHM6y5rUwaDVaodmddV/6Z7pfRSJeDcCWdT11n7wrCFAOh6AomZbVASe/6jmMsJylvdWBuBu
00CnimvuNxoBlsuzUmsOSOgcGcqD4eUZ0VQ2b19pI3w2vGj9vkzl8NLKAegbaii/BydQidJg3Bbo
/nyey47qIshfoXhGIPUNsdMwbN5oTUB1jf/aetTUlauNhCf43riJkfBJBjyJxiiHz3k4muYAZhty
QaR1oynjCTnXB4bBqPuB4fDRfjCfLKQBAYL4e+9WMZQYqhy4BlW8aLhXyK1fs4oOZyFzF2VGZxTp
12rKl7xwRdW3xATcnwQ+McBhOB/GJocLP8lAbqy6vuQbd+0zkH9/CEW4JX6F8/1B8TtO0QL2/EjZ
NlswQETSloiZoMBl7QUcYgfmh4gmWsATxvcsa7swEeXOHlxJ+S2syTxMbfkeTVfWJ0FIVotF0e+C
PTKVHabtFt0ljJF7ndUz/+nQoKsACDPHPHuuqEHARy/+B8KJkaxbfPPAgrA8T+DP8Pc2x0xaX/q7
c2uS+0sDaJqwdifcM/tpFB2EYD3UScufpDcq4f46U/G+seFURxaVo+pbfSzHiLtig2uex2a57VKo
3MBGTvjalggqY9wd4+JvTeLikjkPxrBHLtMjt8CL++bJrcIt7uJsvMhqnnobWH/o29EGD5OQ1e+Z
0WlotC6sxj4DJiZwX0y89iLM2vAePcI3kqqd1auLFgMTehuWKeN3keQJMHPxGSlj6y3FjjTakTq4
hIckBxuHU0x+jw+3kbqL6S2trMOVEJmDY41ySo7sgFGcuQqKqVIUpMvQT+mh6hYPbui6BvqZrNc/
FIEvqq17dH50nN9LQSBV/vViAhwwvxt3LiQ/Vx9feb8wkHkuuvF7+iuC1IWihBAGKALdbDt8kL3S
UAFz1xUv5qCGVeGG8KPBM9LgXXGiycpJf12Ht4wryv3mudi1nScgJCB2xdpwcNBdCHat6eMCBv9A
bbB/TYv0i/d43KBfI4eQcbYEdGexgIlcRuIuMdPSL7CVkFog9sBWzH7TcyWVCpPwdg7JxkxNaCQL
uHlplpsDFkc4/8zSrZEE6kcwje3UhnvYy9SsHyFoF5jU1r9xq2mtMlPGZ95RFiC7aXCKoFrviFN2
HIhAgCfz5CnYwZwowSemr7pGCnqnzJhyj3f6ElhTAvLnNNUkYOy8wIPwtH8mWxOXcmsLw+jsD530
afBx5/+0qhts0wJX+9+y5A4Jf7Gpmnhqyvk2lDeA8hPPz4C41Ezt0BBJNVQUWFWHpyhoiTBLWHMS
Q1Ga/PzNi5SyeRZ56l6+E21dPtOweINCbWlUjDyfLlSp2ndfVKrZqlwmAbv5lA0dnhLvv/DSx25h
zGvRJ2o+Z/oouZCddear+zAjWORJLglYCsFQQvICZ+j0c4EANaUZf60yJt9fnYTyM5ND3K3UidXM
PTpHeWow1YLlxGehh9UiERxBO1czOcTg8h14j7+06xNMmIy1ee73bJ3ZH5NX1k0NRlGuZW5wSHdO
PF2huN/P3f+RzV0HfJUFGDQ+T2DUou6F5Dn28a1I2Yk9VNVIRTF2SK5h9A1sJiexysiwIIUPXlmS
Kg/g7EPLTyeroyl2p58aotBTOuEhsgQBmDgurJ2RdAPPRwUEQkWseNmYvjMxYaOEqEa1xDiytDVc
0pZKRiTXzzsxI/q+EuAUqlmM7ftUU09hDVnMEvye9W3luBsX6foebzo6q7qfTF+5V6b4AVTCzBhd
DAZ+VLhQrVr6rqd66rOuGu3gU1XIULR/ONecEjVlQg1LYI93NfqjKu1X8kxmdfly/jawOpxw2CUV
8ix84/p7M2X8/GihwG0UuRA2TPz4anKH5X9sV2hr32/PeXRT/cZGTarsQX7r1I3aFsa0/+IQ8QvP
cfeJeCyt7bwSbTHAY72rWHUWynAOg+llrjzavRcfrr12z/Us94LYJT8ENZZVkrIYJZeXVl/G60QK
bTVgeAdcBlU6vEbfUWj/KC4ZGlPG/a0CDToWXEuMJTMTOF8bRzZ/MehNt2CpTuEH6dm9PWhx7o0L
8OpCrbRc7jjuMnt72/EbvEJaqZYyKBIEx4u3du/dNKRXWqwXheHhN3Dgg2bVvSNTajX4VCQGSHrl
2KQIe/Cujooz/V8hVz+7urGsySDdInhSzYmEet00qgeEQKCdm9WtxdLI3F5gWb/wL+Moozax2DhW
70Zn5ZfVOLxx/ZTltYwEZa/GEsEUJQJOyJ1C7M8clUBsQV6/P/ACLvWi8JJ+Q8kS7TAU4J5wLK4y
u1k+gTgHYF1tnlgej+HpKhrthHf60sM60LPYQCtN95DeqFZXkayHIVMKliwP28mIR9dnKYn/OxvB
BdZKGOPEq6m8zx0lLPzJZsN/2heQt/VwQjW4qB0sIte7fDk4quIkMS0+nf+fXVvUgMB1ReZFA/A/
dpz/S3jiH5AHQQc32rGIvvQLkv3jlQh/YoqrBkfQhZF6GZY84iqMut9GJ0pBsvA1mD3rU6LUFfDB
yF0agoVNzySGkIkfA5ooMF8AUCGFEMMIVKK8XtkDW4b/0ftdbm4WMGW7VD5Cx06kUkJOJRNEBgZp
0GMLqkx2jaReyhdBC9JQk0DMx95SLNT+Dp92ZC7ljhxtDvjrsoiQSd8am2PhnS+l++iTCZ8Ufp1G
vM9Dht65MkbV+YAL9HVUA959Y2oQ+somNdTYnlERjGepxxcBdxodyTsA1WHbTLR5EKkSOacgyHTD
k6s8k/ro+5GoQpfNGaxXwcLCFNLwvx/4CHkPNvSo8eh1VUdb/pDqEOGguvnB8IGkeJmFAmHU4Rg4
WbO4ko2C03h4MAF7klQG1YRZjNElPEMRjT+V1f+Yof9wlqk4icHIc/tTfuuab6ZLQRtG/QmpoYHA
VXLDsLRpJDxglrTkftDMXGKzUJKEK7RbwTy5GAS0eYcxs5JwVHzH0KGJZ573Rea190/k4mdH6aY/
025VI6+2SRToKrSBhCUvRIhm+5knT7lYAT48D2mTSYncC1irXPW9EeXz+Lmima+tlbtorARf/2S6
VuCD9mGoETRScpJPC9JGMnq1Qsz5dwsae1YWdySJd3572pPP652L/S8ve3/CXHZfEK7AwuKpqnWy
qw17jjc1Pi2DKkv+psaotkAd1BwHat2elNzIqB5laYb+3RDhUs27xrGEowUeEh/aD4WMDuIzwii5
56AEh4C+j1xCGFcgqTi2/PU1v33Z5/WrrZH+1Ri/WN80MlqOhu1+4ab/yDSYRrZZqe6iKlwr0l/H
/9assrq2YCMcFDhhi9DLY0ehCKhvp8kTsb6s55T7+n1ukofdZYfjY+wZiunuWYqeX2j5WwaZoUDz
X4Nfq+B+PfhZwwhVE9nuHdvG3qkY7+a24lhDYmvAdm1cJJ8t5dxHRLXsHEkQJPGd3Ced8MAGJ061
XCh++n0SjIbo25jWam8PQnipA30m+eRY4+W/0OJiYQxBRMV8wRwxH8psPDytuj4JzprX0NWXzUmz
QuNbVQwYPZfyq7hqHtqqJeI1LDW3cQlDeOID45kzutfvgj2KjG/mj1/bLE1bWb03d8rjb567iFYl
n5i5u2OwKg418DxcrcnJQLW65TEWsV14l72dN8m9FRtO8uVomFkJiGvs2U4Lb6xTjrwcysn6ewGM
E6IbwT0Vj4FbaJG9p/JKxh2m6/fmmgcpVv419ENMp3clKg/jsoP44iUgN7wbENry0+2W6YQstK0b
+3v0Z63J8iMlSuL2TaU8bD8OktUpM1CprS6aMjyHR09mWaE3XRgQ1IQ3OG/dz4IKSSYIi3+S1ucu
99ta3xpF8pSOz9kw292AY9ad/vHRNOUMBGlU1U89VOyApnbMbaPHb7UlhOnNlZt6vpxb+OET6ows
2xHMRPTin881725H3TxwOTCs2dp1dQMGDsF4usDx83AqKAdY8n8k/h7z5b6N/y56ybBv4Jz0flip
5GacUoksuleOulax1JM3clUJJ8Hz8kb/c1cqfwrSbEpsnxOcmuJnp/yPydvb0RfDVhCqOBD7MWYN
hTw3kydl0/MPn45YNEWiVDRMVfvCe1R5DIZ5z+l0PA4BrbBsxbHu7bRLk/PzDGTPQEuuhIdDF2xl
/3h2Ih1NNg3CjOz9zIaY5xRTMIyjirE+e5z8Qb+4JUPH0wSfojsTbp5SmVvZkfbRQX7vgg+Z87cX
HxwI1MekXq1XjI8LNJ0eEBrjvtLbPZzZGW5AsYx33mKGVy1Jy8E9+4rWnbgh0+1YJjCvrZ8r5K8S
ggHXsHggHJbjHvFqWuvquG9AgivY9CFVj72+SSVTGurlW/uQF7PUk6afTSRZHhnh/rdYNDAi/LPR
Ep4wAgLwQkH4Y3mLcxey+MIFRAIh9TTiZATDGTU4jnnP4H9yqZdaqu9S7pCQIbcZzZHmHIP8Mj1j
mNJO/N0RUGnly04EycxviSnKYTJfQ0+GbpzmsrbbrwGjOM/amREDs3qEfKLk6sjljgPFjM8Xp7iH
h1oA7So5oaI+rQBdv/3eoFPQcAFub8QbO5Z+bAuLMiDzjzUNyc4yiH6yQYKDnEzR49uwCf45iSTm
HFd+L8UnAGBz3g4Y3z6cMw5bpwV05vAwVOb2bsNRnuhiHOkKLTbdkmTpcPOiID9dyYuNEIlb1rhg
e3ZtRm4tmy2JvvEcKDAbby+kfQ1eV8oQiYHjcNBpkweDz7FbFFRnt5eIpPQ+OFdNsM66QA4X0HJS
0NWk3ahR5KCe8GuiKBfKVU9TTKGryXNnRS2f8q9i+pFS3jcf8c53vtEifv6w8enw/9GWinlAw2Xa
2jws8I2DF0BYsGDpuUAVpMCp/7liIz4qJeNi1eaOEuiG2VR4HPMEMzl8Of8UCvI2Gy4SUEsllAO1
xBQRBpOqFlY0I0ZaAQNht9OIwd3CFU5TXCQqOr5STDxA3fa1/wDpRmuh39f8DE7WvAkaR/ILDrYK
m49f5zBGIXGJm0MqGUyt+aXmBeA8tGxyj/Hva1O3Zs8PFuA+d6fKEDnzmKFWL55VMUf6H7OiECYf
MpJUIUfdL17igrr0UEeuzLfpI3HfsJAsfq5IDbyKTCYNI5gM0aI0cBP9kodAkeiX8aU3V+GlEPGX
VwhvIQctVLMOfJi+D+lH47c2QzrMZX7b6SgzPYioOfXenResvQPFDZviWfc/Zaw+QLU7d92nJ8go
3O25f4KAdq+keorjKRcqAGpL1YqfJLmK6hQxMZAyAU+xh9gxjftkxnYkzFwKQKD9cV68ktR+ePwM
aYAn38p4WYZVnzIhA27EDRCA1OURdXsu2ZuqfyjFJJ6+Rj2JCa3xfh2o0REkIqj5+ykp7V9ms6rT
SF00rgsQhoNXhdl3aDosaY8REMi5huyr59HfIx2Dt8L9MPiAagEAqI3f0h6fERrn3zQ08sxY9LcX
YkOckaiZNAt7N8QqOOSmvIrrv9Hk4TLF/SF8WTxTET9oiM13ZEcQgVDbJcBTgA/CYIFEe5/uNhkF
EAxkQu4Q5gDh3iHm0GMfd3v6XfXIDHPIXAnw4zGLjTUSmZAn+OjtDR/wJzN8fEsv8FLwtdCcPMW0
qWmN2SBwAZXvEOv6hI8Rtqws4y9e08KX7bSIdTu3ygUyZDo0pxx2pLHCS1gIveGuTO6d1AnBb0hC
zTydT8kSa6cUHcRLrDA3Ngpml2eAgS6ENd+cvmAD49ef+PmAKs8hn+hfWHZ+Q5kr08t5tNY9kyyx
wYE3pWJgrQcSjqXEXzDJ4MYvTssFyrLrCUk0l9FlYVH0GiHdLkbcBKuWNhG8tUfTjGgsCYNMBHXK
gsBpMyrOVf4y95I2oXN98YrtqEStzeuSg1MIlFLdK1k7IwpQg8tANoSXpZtGxlB01/TGl3fqm5mb
d7PjD1ueF5MC/h7ceAmpF2+nizdGrgP+Crqs24NB9QymUTnBvz389/ILnaUCq4tpJIzBbHqWjJSq
saCt5Ou3dMeuZAgf7ymmF2Dnj2wqmDVUBAP1pzOgwi1XpptvKmX9ijCK4jHHhzK7CSufnqZr5LXx
OHSWHB8lu8EZMfTN9z0zvh/rbTy3Eaj60atpphP0lssotwi59DmqLJ/vCR9xQdD5NIVpSK6i0o+d
3H8cDyt/gn2r37IOoAHl3VfbWTltdTbPGYkXeCZv9xlT5cNr5tNIwxK91hqKfeVW0h/I2nmUixQ1
UB8jCsiHjZFMphgQCYi16qUUgLcc+eJY5wHYyR+gqwAXDW+Ab6E105Cs33OHIDRRsxnaamT2allc
qpAwniECr1u/+mGDaNu1h0XcFowxz8eMFbTG30jA/vr489nz04JHfvV6sTNXdNJe7aEEBAfajsoS
weYrHuLAOxfxaUKwo+yRvwa72SxA114iryx23ZRev+6jchCf0530nTVLRuDhGHv1vCTFt6z+FOlh
WWaonx1LgVUbz7iU7XawYdikBnWuQRnn6WCsw9UywzP8QRpl7eOntXM/D9ZNcmzn3NSM3SyV37wp
XE/EXETcbQkfxXvOwJbqbGQGGmdjfNke+UCdY64TO+eZpQmEa3aI/kAwP4Xp2YiVI5D8jOskjtbq
ZjDl6DEQHXs3Mq/PsBtStuUazyuiyrfW/QNpOvDkMALFlncpqphbfyt0xGWsUggYsJeUnGko3eKQ
KFswYOrHA0E7dLBq2Hu/A+FsLYa3oNzeatcENMHqYfNduQezap7iK6GLG5a5enAwYiwA+fqGaiXy
hutU4VjJ/oilpNxH99xmjFSK20ni+siMLWfsD7podqr/jXAlFb3IMSzJ1Szi4O7GazElr9nCVps2
HZqAgpkxlv9dOs4Gr64drHYqG19bYL6zS1hOiGrcTnDM/GwGTj8uiYyLfQfZ9edJtaeBOL1zsLin
wDManhUd5KkhJ/ccsjnAxjzGgXyiO7bWmwuUIV7Z9MhXboCPxKPEJFif1hpmCemdayKPeHnVwI4D
0ku9010UlaoWWauqSHoUCtNa3qTct4WeAUIeYJtVk0U+lFGnJQlNA7Cv+d6hmfoyoilVl9jtiZRr
2Db9ICJfRs/Rf2kCgb2bsNPUuexZRNJlpgqjNqDInxfqoTSwzbQXCB0Z5YBO+ExPMhg5frFnfk5S
D/KF4gzHoGdk6RnSb9y4rACCXoQ1CBHet6c0NvFexTSR/1I/0cN9xG5L+1rdQ6u68hfHCeurwTZR
DT++IL2rSdsYBcCcQjVf2esHpyfpKkovmKdgycw0ffYBccNYztyH6D8xv5kJC8zP0fks1EkoN03r
l7P7zgCh4DCHjUe2EYKxgqk5gWUyN7KSN1EYCmJZ++3plGi6WluSTgqs6IHUxoMO7Lo22mq+kbjL
oSQBHOmgOVkgnGuLo1qn7FSJBTJb8rD2JuWAJcc7QxBCsj+XmWjoXdhMWk0FvTNrsLJvwmklsvOx
2xHEVEgbNvc2erylFnrzZOSURO3nSZoMr/r9DNuWYMIqDBf/90BLSrVVZomDA6m3W2SMfgW9gesJ
Dyj1IvElUGvPsKFsKbLh/UByTi12yPNHBD5FFpy4bSDu7mtepAcAZMB5rC6yS47tvDsuMNO0g1uw
AqnVCNaKmW6QhXXoAGBh/quvbmAtZtj7rKTUj0ZLLVC6msOLmsOr4RnCzBG1B9nNBgEi2oIiTLT4
uJIB5BJXUs5xQ568sjkbpUqv2p3n0OlVJA1J+g65ZDaMVTatXlIOjEG4OrPNnMzZ98cvRy77oneQ
plIqI5qmjyZSd7ijddNushkaWZkZUomFroJEP2n0gBousK0MNoxiNu9Jjn/IdS7H99qUwt80Egxd
mvZOqW/09dMpx5S+Szd3p+pixDzr9T0XHqb4yRwUI6LbY/GjcA9AKOtc7KOS38Jl2UszeUPEFv3E
+2T0G7fcgurf8hGxiim64s2tBC0ApJs3tibwKImV892z4GZcVhC5WxMgWrD7dZjvdLB0dCl2Z2zn
flEy+TR5Y+rWEzQTW0kIyVDwjYT5IVsFX6wUQqrCRuQjy6WwnJUw4V8B+zlEU0OTPOYko/LYWLUd
JOH6IxkX0VtbAe4XLYOiiiRWkGhJ5mgtNg1aYYyLH1ewXY5qWHpEkWjnRU+YpQkS5/30jqZDR5yw
OaxBD2GFDO7fVOPlLzGtY0jLQ7r6eVqE6beB+/RHkbB6mamv73iD+6jaA7yoMXmzWigKtH33T79n
xH7l1w+w6iaTHs94olagkqADqrmOH71crNlx05obqzgj7QruD7ugOLmmUmro3oYy1bvn0a0GldrP
1o0uOL0/W7ksogskGAfT3r0zspm8XutO65U6gIgmSY4YQLpfk3umiR8xKD9/fEZNX+FY7f/I/qzA
V05USGXYxo98HoY9iYGwjCKnd1eijkoW1oHxPohgR9UbL1hAEyOmMlW+oy/lQ6/EnGoZVzApOlTR
U9jhM7tyqNBKmXgID1tpMJpLq55XGPZ5OK/Ef676q2ORQ0kqqeB/0rfH+C0HLjmOXb9yiQuBsVgP
TW226e2zTAVf7JhdniT13mKqUnfDiGplur85Mxsjpf8VmXGbg5GZOlFmCcoJy/0LTbLH21Yemjg2
v2ae6oRVYNLSFH8nSsqrxu6+vchnwiuV65bWAQ4C5PxvXbkN7FCGXeZWWMEu/7mhMQ2mKIXjgRev
YRWDFTZjA5ilTVPKccT/JycXkzXrx2FhvX26w6NC4dB70+YlgvbUu+fesUbfPi2F+jDYlo0JHtb2
U7+YVqRv5VVQj/veD0t0MO6WBxU9TGYbFobyw4Zbh9WTBXN1LoKrc/e/m/gYTIm5TFoxTFYeVoh2
ntwlNvToRB/k7kJV32lwFz3zeFLIjzsLKAlMJ9QSncd3CrFqbciIltNzkGvrtYDq2IvNLdC/8ZW8
vi7bMGfi7ZK2I8a9bSImnMjFnay1p/Nfv3Iwliiwp2rpNDGMYM3rHMJE+8svGEbvXyrmTzvxgECK
KftvPVPa9prC/Wkm0XHEOVfyNLFLhxbPeBgJO/RdCEPnqc6NaqR4fUp3uPQYy2xNA6PaXQIYHbZ5
FD3rC32aINl3uPOsr9R35JfpQ05SP6NLWgokI3msPxwtsPSPJxlbeSHT4to2k6FfpUbxwvE6fxma
Pu4iLEJVxfK5LvjiSxYyv+HncmcTMLKp6sutr3onZ9+EPGJzbNWYVAAOOXZzhR3aqlX5/l9BRYPp
pwsJ6NUXXRhWfPi/d4SLgznMiztWnAek6Z1Vk5cYnhjZkl3tfxZ99hGObG2KqvWkTGN4d2Tjx5QH
kPXbwjjD8CPkJ5YL4lDlJgDeQEiZ4kNHBu8/V4DuwsG1z0tiOsj63mU3puGklJ5E2tsot4N4gYeR
W9WnJ0yW6XkMACqJc/fbfab2x4qC5HDGfwqROFqgP/kxvoj8P4VoFvS/bYBwztdvu8zfy1vV0tD/
DG9Vuda4aNzu6ClDg0yrxEhCGj2g5GEc4dv4R6aBx28c7AMv3Bv2p3u7RborNOvTjeL0xNGvnRdB
tdWuWo7vi8feZLl4MxzAno+hgnN3lNXtVJZM6rk2dtD1Hm4eM9G7jZzy9sTg+PzB5SwerQjRl4kg
+wxisD5jNP+NTS1HxUp+U/ibyQ44483ZucMouY7zYZp4MMTS89JarnWw+JLIBoFrerzxXWV64NnJ
oBS6NU1bhVC7iAhXG3bgWPGrlwpllkIk4bl1VhI5IN2FRZpnhxFUaVqxrHqzQY3uqaTGFjs8H9Mj
cFDUm5J0FaXsXI4R0uhVpA0VTXz3R0HKhJozaruZguHCCHfUKqe0Norj18xKBpl8YCCgpngZWhNq
d6tCgzX7JdeniBjNO/26Muw6B6ZvrBRVOdViFGlOCNEP9jkmo+rMN2L+MoMnHW+kOcDJirxswxps
zjMbWZs9cNnLDPf+0QEqMYJ+55NkxrW0eHprSQeh4744fJkId+LPNBGrUKLhTuD+jLoWaw3I2mGD
FjFaKc619HopLwzqacHwlFxG14Usa2XHZIPnnrglbzkzzT8LQFoemOItSfac0EH2doQKhj1IqNtl
D9U9yzhjCW+/pvfO6dmZOtvBsKgWLmDA63LOJeXQZ25InA2rKl1zT3gVG3G4PWOIUM5GbEDvl2Db
3r4vuFMcAzWkOAEewMK+blO3qF+3rJaoH90cLmshTGj149RCvDehO7+HPlhVShCSlaR4j8R+cMBt
qFQVAyN05VCskdxge8fsU54xyEk5vXXihAbHDSMfolHeLv/xr8HKIj9u3UfMFldp8N9PXFrTk+ZS
/qVdW/cOoh91F2btBdOLn/HjMFUsuRhZSrEPPe8Y9PIr0/LAvnw7IC/oT7OaBIixGjamGG4AAC9u
NgKJ/6FgWiW3cz7Qic0rxMxyP1esmyIIoz8PmoMBRCEIuoeH0DOpqhgzQvMK/rDuv7+7nWFGLiM7
el6PcZFS8HXYl1wnxe5kswva+ZXUEINqDqtkRVX8sMUbEdUvh1a54XWx0UyMq4O3H+0+T0PSdRmI
JxYxWeGTcVt+UZ9ou+ACUJDypCodoqTG+53ExIdlSZhcaOMtuqQAziuPp0G8rVLUWYXodujuA/Rf
tJLZkmEbBbxneJKvZ497NxcuhIZoIO/SPgHgjAtOEqGa+JRoF02cKmlnSXT/H9EzVjYkxR0tP7hW
bGFgSaGuXyRr5EnaS8mY2N6AaEfwRCrF8o1mWsVKBzWh4l6YIrVy7mwxM4oTFsX8XxJMfSQovxig
+ke7w1C2ZoKbfyKUjAG8wCGEXGP6GejNnCr0yxRcC7lkf5DiPySeFbCxwqLXV0ffOi7PEDL/5i1r
cqk7xSYCCrGDkBOZqAEF7LJPqBMl1z8wMqjZhNP/9ylrSSigVFKF1xdVApXpqDwnqzW7y3kRilW1
aTP8j16CLtTlENgma8nb/glHuKkMboUlbBEelJnGRDb1LYcFKz+E7YaLzCWnOF63/2sArWQo55CV
pl0gaxv3P3pZ6hvZ1RgwAmDfd6KVVciZomr+gYwFIW9rNKfyZCGrC1+JU6Se8H+7Bfzo+Ozl826E
OPRxcyKBnybYEn+tgfwIH1BAX5mHPQL7zzgDYug5Oh1QzZsrrLoo3KgQZnhSdNJlFzGGK0aPOyI9
on16tq5frBe2oTLpuvUleKGMYc/OAM3/rs4nmEbZQO6avtbM83l33JfgdSQVgmzn+TsE6LkzN0Ym
lGKsjWEqaaRcoY4JQSha5puboMqLJpgzhFE3i8hPs5AofGUcyp6+OZQLsGJ86KSRT545CQNQS5OS
BPr60h2cme2cRwQcJKa0x9wjJQHtF3xGloDN3GoVjcM4IjwV+plBUorRb2c7CWAv4cZWEoy23cjK
OoHfDsLFcyYESbwO3t93qMbmiOfkUhcxNWggk24V+iStMrj+JKh9nkCuxwgQXQu3baffvYF+Xx8A
4+0AazO3+98gJj4OzMKEGycKHj6QVsG6iZ3zpZtRrtDgG5vcYnYKLx/t/Cu2UrG5+UucrmFhAA/7
xsgoL4QAzk+QxD7hxnM5vkGZYJehC7SFpPAywxtYpNqXRgWwAk8SVovKZ5alr8kfpQfM7FAmECma
mzPjSXT1TvphVGxG8FJEtZysNr/i6QwybtpjFlQaJh/IeDxmNusNuiLCkA7vuqurjQRRs+25tuO2
mG3GFKrFU9m9gxv1Pu4ee9W6qs6wksTIh4KBe7DAaC6qIWvl6zygSNT5AfYZKcMWo1+fWb0QNBpw
camnaCdhERoGBW8sJ6e6xtzoUUeIphNb226sHu3CzK2Phd3Qhxk9o+jHLXWT8UeaZc302f4ReuL5
oYoX8HBQFcMpHp5BwU8s3NKqkzKYXoAPk5OSEPwi40f0+5pxSQPsf3km2fvAjLaLvFeupDsBNins
7tnntn1NfnVuqxhkgchXLideTz+FMEKs8etQSNqRxbICZaieoe/rJwg/18/5D9JWdPQtTXjfpEGk
cc9nOEAsUyldOOmv3w7fdp1wFFhIDStHb7fd145AjnRFun4oFSD2p0RrKYPsHUEfFa5D9mtIKjgl
d3bXn5R5MoA8KbVV2BXeZ9uS47ndLDNvfbMf2Dr01nLqiB9v1b1Y9fon2btiwgHCjvXE1rg/IevD
ORC9hIdIVZLL80tsdULtAmdEt+Fgv3j+uj7AIrKwVg2sUvVDNmVJPiGSEpsRiiM2eOUlaS5rFgPl
NJivrfbFbqdXJELTfs3KOqrw66pFnyrrCn8Mf1zbIWDsXLNAvrfuSBsVlSWpDALcjhiW+KppEwtC
i8KngjaDRVDAR15etyeKSl50xMZdtAiO4S1q9FBVJxU6w3pT5AnnYbTRhobqLKF2tmpWBFPi9TxP
rT1LpE9YPVaR9FGF219h7JlzswvTCVbFHQ6NLk8VtTMSQcpfHYWWPuWf1Nl8rogxP1OvFUC+UMZr
NvjlyKespI/1NL2uXe4rnh0X8+e754guHMkyk+GdqMAN0nQXTu5SmUMyC6aew9W8QPV2viTyjfzU
3ZPV32RlKIimZMCeGwJd4In2KIDYhrce3NcrWvIcT20hl3lG9Hb9sSDd52cXcGHaOFfB5/2/+lFU
+gVBHF+N2RHFIM8VigbSV/ffLbqD1nJaogBFPhHvJpZ1up0e2LeX4KhJBD6AGh4d9UKZ9LdYkIiE
31m+ZiSO0iGYwsao5RZJrzFKdScdJNKxHDmVdR8Wlm1UgNMNTuIGg1Uo05Ja0b8FI1YjPVF42Z+l
niNxFiE+WBudWDWRHsqOtrXEAkG7FRpddyOwpzfaY+0f5LGT3LSdgGJLInUNDKdQjFZRaBm0O38k
muyShUfaPxdgasS0gqwBE+QaIzVAQKniUoazs0KWLh3Z29SN4maNuF1bF98AkttwqFmK4sDVRkB9
+mn1U1ADToi/5/7D2iOYt+/xW+0HcR2v/KxVxZIgRkJPX+2qBjnpr7z0u2Z58MYckDQNGLAimUyb
ZnHy9VvAYfa7+Zk/2f8LjD32xLleBNL3g3kZ00Vl4PNDF8HDs8Bkc1mlgI13o/jzNRloXw6DKxOs
MmhhhLzeIcibu2IwYrgeTSwxEppvRYwxM3PC3pQYiAt7Mx/Hk2RaybgqCYBjRrriyxdUjYrtwdRy
+XxnBhOCbSiTgGIE20f8PAeRWPP+czA97rkFNNIcM5ZeB7yJs/6jVVWL+J5Rj7XADMD2VZvdCVvu
AH8QHfFCWbYR011hSuTujoYxLTtwUm7ttRsNdJ3KfyB4rO+UeCaTviy+7OQy9lQbTnDKPToaS1zE
Ij1WE5EMxI1OgWkVVfKsDNzAIFKHAZ3CZYmZ3bft6cpwgUZ2SLjVPjsykhQeV/8ZV7Y8iNb9Grug
ZwLHRH7MrUA+YPE9t3epTWhyIE6//8xvAwKDqhxhMY02iS3j5YBGaTaU8W1DjqEEsIWlX//7r24h
cLWYtnoGxiQWOHpv95LGX3hMMEEFYlW6HWPCT3yh+bYxwvw/VP6iS+nb/XsrpoTBhQv3QDxyzvQW
20xqIjL3UOgjkrYEFYOWfDHLdFq4ocHExA0VJZzTk6VHcnm494XigycXosS0AzNgGzGdWdFoU4tJ
cMZJAo3Lybmy0EdBIc3/oHBmxUzWgcFEyPJnVFWlPMEDm9UmzXv221EabI3yLdHWz5UwrOv5KvOh
cGevtg0QLBPU784RQP7hcfstCIoYX5VHV/dcBPIC83Fu0XRb4IlISt7oN0KrOD1hcKHgvUHOjoVb
OP3L2lSI0st+iqzKlaD1uHd5qR6CFOhi7FzJ55nY8c1kaJZJA4VA23Qn4zFM/iqXK+YpS3X6SJ08
8xRSrNMFLlasLqJ1dYNCFSm5U0UNqGhqPQn4LYKtIxGe2q1bjJP7wjODRUaVrdk0ukdxU8T+S/Ra
I6Sjp4jjDMMNXLlsF5JKnmvLa4euk3wbjCH59/gs5SpwjVnNKh2khgUw7Th6Exx3vKfqlAjuJNDq
fGe4TkXMFQuxHHeOGxIPcV1RWkwPEvlF4mWZ/vrxTSOAN27H0sa3UvcXFOQRiKTFGafwt53WTHVw
mxDqpQgD3dbex5Ii4XZNL/ni5G2kIAuxFVyqwYbZHUUIi9Xi2ngQzYqdLJYU7tPP19sVY47HiqKT
dOPGKmX9eeWWYnSFWYo+lJhsX2zdthMuACP9troYEqCZq5SdmtkFKp11/kRHhVpfH6e4AoZ2B4sC
YxP8HDbRFxUEHFhZq8sjldnpiX3CMA8aTqIH1X7fua4Bq8OHaC/mqUlVGuaGKFWDiVtMg6BxuAvG
4aI5IygVL8taHTvde/8S9jkBW8WSfGcLKHtpXWRFj82xZ2trW4tOFTiSDibORDhdwt5HvoowlOd/
ASeczRYcdlEHiQXfjMWJXHkvi1MbdYj7B9GcksE48R7mejKLR1VuVJxsj68WobTwB1y1RZvmyyv1
1GKJnRkq9BiGA82PBP9WWB389/NhZF6Rmn3nKYwt996T9GK2ERWOdVs/mh9sTGI2NmBgf0cFtCrA
+RFr6ZLlpIDGagwIRVHjbA5o0tjrFn5qrCdIyLxSfn/JXeYDndWZ4saMbNZ6J8Wv3/kwsv4EV1Ma
NkaGEzLPJLfLrTB5u4qTOVO+kSm6PC+Xil2Z44Zytlx0kQ/NxOC2CnolYAIg6B6eThPLxJsBsDO2
F8aTkoF1j3nMmXCn3pjQr9ymhi9PZ8d3xmETQrzNuc1hMiM8rK8Ql81r5P7iABP1/m4qX5F8piYy
qm2peBANl5SJn6JYqrGlL7B0F8zoJNXZaGWL+gdNvhQeK8cscWEpmZQr2wcIBGGVdWcZOA2KjtiE
+iJWvvYLN/8AqlUY2ZZevKM0b1Xysis16cvSz3sZ1PyL8WIdeGEjUe9/clw+jNnkwIhHjdu72Sf9
H2Jq7C7uMbbh7ra0HM/jXPIqzX82lJcfgNHYrkiXEBiDO8GdnuJFwm6ZmySuFTszSnVxRb3jRarz
KbAytoTQwGK8mHkJFODaTH0lNuT4v+BVTOL5mdoHfY4oNLP/P0BEebgPQe/WK+/tGhB2TtH45vcT
wnj0baTcZhxU242raF9I1Zy9SZQVzMN+x8oGqjOR8aPbVMW0YliDbQkKM71U4QlMrZilw2diwv/b
S5b7mMwfDre/50lEdK2c8o0/tyUvCEP9qIj6cd/wBWeFSSVtqGhabij12KPorI80PDRm/9RndZhO
WWVgmqqfQs2hUxG7s2OFR/FFy/r78KPrlg7+zGUFtiqCLdfflIH55QdrkabZoRpR89tudUY3zxou
hAzl/G0fdC3cBzf1ceRK8EzWA/547Sp7ej/2xFzRWxjZKGMf6VPvPh6CXfCTMHY7+Pjl5YFYOQ+b
aDYTviHAY05Yr/peZL7hkkFQcPd+8fVIcrZPxRH+9L/5tbIfbzWxEomTCAu8ZVUP7TyLb0ZREtnN
5OuOoxf7Yniy/XXI5rcm80KgLnjEQaX2jI+D8XS4TXHxNmUIPSzC+gGK+b/mz9QtbnaTPWqSdxUw
Kk/5VVBgdwjKMcueL9QZkWfwBfjNg8VW3aHuM+M3IEdykRzPtlCALBtWh7mM2DqPP/uGQsO16Qda
wlU1M4301wfvj3FJUHrLZKSH+kOkRTbqi+KjBKKZayrMyxaeQnB/qi67bnF9N0Uvpqh2akY3gCqU
W2fnFPw0UGkXs6omYtUtSNMcil7QZp2zQE8qZ0OCoYuCxv13gLrCM+KsH2ZybWW9FhepSSpUppTE
f4CcoBS1VSCMApIRQMHhqn1kPVGrRxN5I1KG+rdfhW93GdTj8Vfhz+odl0SNI4h66oWQdk2nRhuq
rAfn7poz8UPF9jzXMU4N6TOpcuRqtETpwLxlMfXF4HwqRchexugs0JMRLgyFOQ8N8VqENTe6d0tC
Jvel7hhBMxdZS4kqkhLhnggI6ddfj3MgEG81TN/zuKI3mjtBWrIgqxJw8VS868CCXNv5+8CP7qOi
2NZ0CnzEonMAVTVHq5gz+KwAYt5NH02kTBjcYTjuJnMs5CxC5oVu4kqbWcS2IYCy8I30FMjFagJb
+44IVgj/WszkxGf7Wsiiw9INUlsSYKf1BQ/oOADCYKAG4a26OpNbzRDm4uthxVlyGogF0BVLEXQD
W8cm4HEt/6ioVEvJQE4XS8z/J8OL+UwVdve+469uQ2+q3VhgEiGUD53zFli01pVwHrMgb2x5w7gj
BIve6oNnkO6Hogc2ElaXDyJg4rk0kpt5Loh2N9f4jjKMaqf2CkoQ6Gx1F/hDKFKAd3VgkYXeBHUr
+7YwP3ea5T5o/oW5vaFyew0/TfoKP55XtP5nBUWtuLDlPVVoE7HMGKQKyjOjEkW+GYFI3IhJNDI+
u21qRahhIDt0MWdiKT8TJLg5azWIB8AsnnZJYTk6xOjS0+80FRarlmdfiuewfEJoPNOCtDxVWtIB
B6wDR+wxMbSXXvhFC6aKdXNPIpRhg7nyV4BAjyKHd5d2Fs9Vaps84kqcA3SbDsHXfCvzCkF1wpeu
3AiIpO9GnMzp7SB4JUnkDUr6IvH1V0f7JWLOkOR3WkG6IA3LAsUFQ0LOUyFBAUJeBCPjbZbKJY7y
GaWBpZVdZa4Dt/WGB9Q6SMAdEz7D1eulSsR+Rfe0pe2BRktrYuO40iVgSTiOq+hkl1AfdCfYsBPw
c9v+5G8i6ZBjbCBd9ANiIgPSch/2VX9FsE5TQrlxQu4Q2iec9WyBSPqbDkcU8bEuw0KDDTwZu3rW
XxfdH4nSyM6Q3zmpMefev3jm1DBbXcIHaJNqlW9MVsh6sNCvmVwFhX6mcHn11soHSpNlZJYvYbfL
q1LbLFazyw2QiZioawaVr4UZ7wVhaoIedLEdt2UUbwb9Vek+VkuV0UHONmQm7iunmYxAy0ElWDKZ
/+Mo64a82Lx7p/QM4k2PDJ1BWUwnzrNFUnJDL3yvYah5D8cv9MW8OYCMkDhpNbL05xtSY21+M5yI
zsYYj/41QxtlLwVILMb90WlNhqAnLgPRPkEgWvqq3UtblIThCe4agBHHC/5z0SROcv1hISeMWJ3j
JfjG74L+UMPty8WoQBun6bz7Hifw52RK/sFG4LvUDo31fWIEMvn/qQNlgRfWHX2HPimmoXifcTMj
5j4gjy1McciH4x2eNicMnnEwQVfHY0KcQxWZCJ66XWdouKbZXMHWaQAoDmxL7mqB69zD8H/2JVuU
uVUYzsmMxdtizw3a2mCXhTIqym/potI7DK+6m9DDQZ6i7SEpzHQw1okkWc95Lqu1vltqBuI5FNkI
aziaZq9VNJprbg6s2pa38+6tL8CNc54yc1IiVl8PFt0VqaCWT/aDaSbLcAeDjPVu3yUA/kBpYf+d
A3ESFTp9YRBiUYWtPY7lFTzwdQA8C3dS0Ug1ehIXnXUCO6imKX67z02S/S0mdEgU4C5+ERX2OAMD
Qnje48eRPCf7z9DQ/BZ8nHIlXcQr1MOMnP/DFsJbsnLDR0WOvtayDBE38UCSeNPrcd+Tk0zhRD04
SRaLvdJJ70/jwgYqMiB+E7aq6H/nhLwDrQHAfxOkiVtBFwC7SlcTkCNgtZWPF3tt2ic0VCVWeAwP
yIxk19SjDFpsLFwBO5udk2DK4sVigT+el4BJhKVbGrHcrNZJZei+X8ci+jqxupMULXOXCLA4lrJl
8jKq3Kx92J5Zq1OSI6W9AqQTaPrkeuUBcAglZpNrm18S6Ikic0aGGNt+vs6B9E/XDvHp0rXTCJ5F
zoV8q8zbTTtR0FuUoEerebRUkenSd7og5aC84CrHre6Gq5KOKXBQHCKDImAAvSB7esYWc76kwD7Z
dOpPI8Vgn2/debSrAenZup1I+/n2GohE3SBwJB1O4g6R9fjb1X0w0qFvn2ZOtrfHZaExFL3JI9gR
wO5b8+D/iUIzthce8WiPP0QZ65JTEi6sa2t5pfdf6F/R1VwekVkGjsP7camaqsiegA3j81eq93wE
sgeMXi/2BEqXbbw9PhAmbIl/F+9pahs38uZVpyo3YcrHQI9BLm8gNNlSA8Og7sPh+k81bfh66ZBz
AQzeic3clGTCcLGh2P7ucNPpW7Krcq3qiDOpDFbgtnyYBhZFYEB8kTmymKJO+gxoorkNvGJJwidZ
W672iwgNYlgQU0YRRTs+L2rwJU5hXU7+TiqYQDhBTq8qY4oSUm//L9q7gz7X/IKwPmNiUsuyHRJr
C20SZVlrZEw2AZ8BF66j+DD3jf4xsWlJbJECmfCyd2kr1ZP5pFrHHWFrjRE9J/RLDt7oNhDF8t+p
dzqeYIOqdYirL8GZkYWKOPMTQHYO2/nJVwiC/8M+QMymIq2CXhUSIINm2U0GvO1al2F1983fug+o
c2f2nMQ4gk1B4qPWBpR7a8vH9cyTCl7I6iG9TzLFzAlNgvwJK8X8sVBiYnrH0dqDBnuzN4R6s5hh
kp4L9i/T6Lh+fC6R7ou0ZutsikOy1KbVkZ2Zo2wN/yFKq5YfYUijY+mPG9QnzgqGZ+TN7fqX5SQF
NgZSZ60azhJQ/pBD0E/HsPzmg2sdTA/WdSBSFDGO3TVyiDQvkYpoBLfZiHwwsBReddBYy183I4Sx
xyxDisC9K83lGeKpr+FlIu4x8eCk8Nw9sRLUhcJwH7FqKqLhEGlLRokoQlTKIO9tpJypeVDDTwT8
GXd9WH6e0tepcM64brbuxxaFC+FgHw+TCfc3CB34VxLK03ibJ+GEUu1M64FNAwTKLBvRyFfAMna/
V07JVfLrAVDl08hbwe9+E0aWEcsuwKcqpysM2Nv59L3j7muU7quaiBNjDVsRgJNDxza/yyAolwH1
K0QW+4693PrLSmuCb+h3N9qO451Cy/oFGgEITq/PxdskKnepg90kRr26S9iJcbTyf5XOv8nXugzC
6evpD6nrwbLxgR28T6pRfSWn9CpU7jZ6RySyBmnbS6gi8Q9FaQ2qQz522yhHGonHP6rTdTnsalx+
2T/5CSC9UrlNxQEyFCrWOQYO732fdCj7sqltxvt3zD+6Fe5gPNU57gdpk89RW6hSllc+1XNe1Wvt
jNwVUAV52+/QkBlQAOMM/BbbbsfKCVDGXWzux6uT7y8s/QkllScWaqZHTxgKczDq3KnLHzI8tmMd
VkOyGt/4EQtqM8uJCU/8h5jiUWb6O1cC4C38OWV3PJhohaQ4AggcpJLqvQ54W6tMpgfTMaG6xKCk
j4AnwiM7x8cKvXdaaZghdM5jqxr6/Vvmb50xuES1PzVrEe+AsPhjcGWOS4ZtyX9+KbFaqPoIv3OO
vXvBjGA3snusIqLPay2XVhgwziwNc4j0oARSG7bv3odB4JPObmnr8m/mw2XMpIvF5W+Hb9Xvb7dw
4QkrKDHjgNr05c+wMZ38o1Ozg5gQ+hOaJFEeiuKY+ctfDrx58mX3asNUgAIziOxeab8V/yg/gj1e
eD0+opBa9JtD+yHQR06RunErNF4izh0xsTZITFjffvYRnOZrBapCftnVu2em4USlhDDoMFbRsZdV
KgLQVbrQEi0og3TFr4Z//4xhJKWP6HZIiz7ikLNph5jp0ThtLXpgUkCyRLN6AIwYkav6UDyCvGTK
ph/MH7nZCSCMqjnDpHj2FQcabEMeSGVpJFw70BT1bnY3ftDxb8wiXzOSjUBoH6ThzXVUFlRylxSw
vXB8GDdMsy7XcngSbKgGjFV9kh8N2Up5nTgviwYMC8O7sNi/cf2FZBOpUsHOui4yV9j3pZnj9dFJ
uFvs3gPmubWDNqyxN+0EQoC4KedEtPg2al4xmwzq7ozoC9srTY6xuWgYnTcQ4c1zDTDFgcTeNHHD
DzfmL0uIXsPI6v2c4tNFOyIeyrYOQJa9aKr/kSNPJylQdrR7sf7k8O+9dsISKzKfL7x6xoMdDRCS
Uv7zIFF+SWz4TMgqCqjxArhBxxy2nwo3Mx5XJdoFYHRqTv8+251kGLEf+c2AicSCjH2Dw8jncH47
P8ztYiSHQz8IAJwC/5s+o8UetBDFjlTlbUkZdfyZPiAi2PRWP6T0YykL0RyXaiWXDwsKbGEbNGWj
lMq5BOImP1agqkmvr8pwfuymTCvuHsASVDmh3iw/L2Mg3tCMXpPilXyswJeg8MxB71tGbTRC+hbT
p6FGVhYD10QQpTouVhUpfS3TbFWWGKJfu9PapoMM0SHIEdHll14Kcng6dmQ6KsbTHyyHurzyoiAp
Iwo2xel9ESVyLkn6xSqhToO/aG8oWdxzxqsjYiUvbekJ2EEJPBkcOES4rMn2plygHohUK+5IXyIj
2D57xM+vuN3GRDQvdKaK1h61Fufsmk3kl4ALEb2QIt49LxlW7Xmbr9aFN4WrIjl9XRu5Iv5TMr/E
OLuHca2HpHFXYUMZ+AjHywDwZ5M0pdOEhGvGPZlhUZc669NCbh0k3/cHQms0CYkbTPiWXgfce/dt
G0cDNXd6aMBHGKKKHHID7/WWPluqGyw9+4uiWCguFmAkxJS3dGegLvyD5QEbZ0+T5NMV1sONTJOu
e0MWVKR07Jx+Ed2Biow5Rz4NsjmYBe7WH3PTSdMEhHj8HSVIh6BeE54XeXWq89XBrVH/2oKE8ii0
tvN1CLq3xIEj2dPkgdRbQ6qwVrQefzr1LslkwppYgtYkKzxusQf62lQuceGa1FXiS/FhynSpucST
gAf+0wC5OJCK6h3t9EWviLz8X7QL+2e80c3+fHmJbPj1p5m/SPOw2LtyVZSVwN+hNguf15odhfSL
c5pfgZMNX+f/2kVIoMmnswzoPEJO+m18z1SPSzX9EPj5zlQn/QwWcteafCTgJvJERLc2NcARi/Fe
PCNDkwH0uHocrnBqd2SY1XI8cBd/wW9ntQ50FH4Z0mbQQmBTehDbeamQQstok+fPZ9bqTy4rhd2p
wBZIzfYwTB7lyxp0M3nmm8uDjZsAe39fOb0A4GcjIZYkJviM34ShP58eiFVP1jXSLPIBFDCQgWe1
ALy61fFo0V72eZXHiUG5SVGV/8z4996+BNVeSdmPsXhxahKWw9b+ck9E/lyAJnDk6++sClxKX+OF
aiUg7Ea01PoBtyn8/ylwcZRshH/s1kI93dQS+9vYIYt4uLkbFxTUKx2cvTwu8fsleVW2HQQ1P2Lk
tODLamzlL8f5dI/BOF0WIC62vG19TwD/c2DqIVtzvQx5uaIkD4hmcVdssaDQnnJa0Mitc2tCz3+e
N6yNeyKf8tKdTOk0voSSCyl4oVSGWKy0tuGu/fPIXrsEELoo1L/4QLC31XAmOcm77+4bYwYqka8e
TIz7sFHJi4zpWyhL/D+z3jiV3H4Wc2eCl5o8XvqkzEqWCOO3lqSYLj6ivFqbt5K6W6dZdND79Pyp
a/n7n2UXPozTcf+ciiOvCVJegCu1+OvNbQie7ZKcqDX8an9mQ0uVEthAfprhl6Wwlkhii86eQ0kj
IE3vEMVCQPEx9MANeoK1ECfu+6hSEWTenFiGe9WbtuXY1cwyI4B5Ze5HBZjcXO/+PsCeul77tiRn
ekbQOg7CzNlq1/w3wDK2nD3QXHfs0SlFXEOmZoXGroBys6djl3mTJa6WpcBZSp99AOLTRUGkYqau
rPsfcee9khw5VeTjf2a+ER/HWdv3qwzyotx78ldC7FjYs3sjKBubJP/tB2aleXfP6RcVKuHFnY+k
OI8gt3ZCpO8vi3BRMAkdx1S/gHmK+7/gzd23rnw6UfiRFz4MyHUnJtuogP5Oq1oqG8S9wvwDnnVr
7+YOAv8Dp99kgwYOjQPFZ2TKoNptxwgaygfu9ExHCC1qXaV1qqM1tdF6aonK73cYMzioBV8PSfwE
vwMTi2v3o7/sg7JDhgnIXC07fdHi7qqqKpCs6KaYUbZ+Rqbv9ahpwNrQ6/lfhpnxE9Nk6Bh0MVaq
lxNgywYsGtu+zJ89MBOehiiAygDeejtanxp0hFZAZjdoLPWeRbLXbPlfAsV8r5jgy48Vfp9Ba2Zc
0hpUO8OxjSx8n62l4zDFk5RwwORCazPaCdP7gZK6gqSGe8OEzfci/bg/RzMDNKHH/IW7JIyH7tFD
Z0lFFaIBnnI/W5X/e8xeEv96hlUkKK4UOo/pmmwyFMmfwC6Th2MXR4NhJk0QuR+3N1SsxOEJ07Zc
cxlMWZsJLugRFE6RSQMNiJ+P8uuZjekey9F0ZrLOFc9IpJRo6vmh9MJ895zh+nofLD/I0noFFE6D
/33/OQacNvu5k80w8yFR+4WRs3uo+YF5TfJdDtFBX8Hfg3wLWW/Vv5GPocAXQaijQokx7fPGOO7J
jH/6dOkq0zSPBRPSOUNe/w6bUNID1eYeDg1njW1+rgDsK8+gyrn+rE5/hp2ILJd/X1gnHy3SPWTf
TEEB9mY1UQ9i61aF0yG7mJqg0vj7gdP+3xlGPimCO5Tj2h5HcDimSBLDScaQKwPSD6jz3Yu8GS7h
Y7CBT7MC61NHa2sWi0KiKA5psVaagTG0L5a2z3Ufr/vkR+ovO5dc1QWa+qPINMIy2n/uT5Yhw+Uc
dFi/CaI9dHLe21eFsVbmtEVCI32lCIhQLSzhKxq8EXDJ/Hf1pqlnRWYwI+dajU4CLjESwdGC54+n
GvcETDEmI3ngj/x8VGgPmCUYYE7Hi6kxJvpF3SR4J6MDqPDenGcAZtl2i6H6pyKAXC5G00fGoyQn
vcxYNqui89mTUd0o429Kc0cWHBX9nsP51h7I77rq1TbtJIFEkBw64JeG5SotSH/uCLoPX8ZQ5QeW
58nHP5cuz/0apaGK2a4awlEQEIZAWiH0jV09KQIwmw7HbS8IfI2b92SvcEwXd83B+sSByklhwSDl
pl38d1MIgOd6vGyPLom7b+m6kpUB1sxNhuOeOfIHGvPRXjGPNeHyd4rRqV8SfR1PFl8Db9bHAKwQ
Ero8MnKju2/cvtXdZDg7mpgvjLAv7FMiwC6cKy4z0y7vqF4ZTbgVEqMHxmSneHXhZQbk68wHVxj4
cuU42iFzTsPdBYzbQ2kdbv+aLCT4VySvET8Ca5LG5Bbxq8N4d7PAgcq2qqUI8v5V+zWuPq3thYPM
C0rH+ZAtS9Dxs3lxVAgVuhQkK3zHC075uZwdntfvr55BcmITLuEkgMdIRYRSl6EaBFV35aBiEXR1
reT1A5YmpbEgNkUgu2DOo7UBs2wKhiKVPJ9GZOdWeCON9mXmuhuEnmC1E4DnjHbZlqTcDTl4qWDN
1hPRlYc1n3jYtX5IaCREI2kYL/xfMzwN464nMrkFpH0hJu15z3Mnzx/csLcjKo1JG6Cky3JkhxS1
eT0xZgIx3QlMB8ddHedWyGUWSKUze1LvchrYojICk6uR8reM8D1IaFasaPAHcE6lJaDVCSoGIglE
wveuef9wpesQ4Oqv5ZaKBn/Gg/CAJPiwM/KyC0I5RhKKcjhzpM9m5VKDrYgtX4tIDYNXRQ8CjqZ+
87uWFdH4lUiyKNGV3m2rXgtl+GLNSQ+Pbxz+V7l1kWpGqvzdsqqK5u5snT6TQ+MkTYRwnEKevfTC
0KcTqPXVR1a98AMUhW8c/l5FF2MHlDAgyrUGe01d3E8hhG1SNcNiWXbC+U8iW8AgFp/NfKJ8gEqc
1YVBMKWVaYBQDLeofBszGgsWo8OD3dQnnaMWCqtLeJuFPMjm9CHGd9g+V0ekEugEspWje6KvSZoa
Ttb1HMoLmMdd75B1dJj5L6chnK8Sx6aKbgkfy3CTYAcOyMmPvl8ejm3yIApHIAayz9IfiKtaDlHd
XkG2IaiEEDRZ6S/ikxKmJvcyrLK3nhpHpPPWZg994HNfV4xEL0t6BH8EawPSEt0DMTEgPBWf8fg1
Pjx7uWHg2De/dPJ3oa6ADY3atEhgn5O5OSY9z5y1xv/rUiV1xgAPmoURd+xRus05rH4YsH9GMPQ0
yeYR5xjJPtPC5hI455Ao9Yxh5hJ7T2qNU3JD3G6vhVHbYcqRd4cvOcWr4XhYW2f/oBvD4Z7rYS65
zI/FU2aP2i1t3rD2s8iL0khcDKcz1osczg6G8DFOC97JuZlEEmIJOpHjLU7G1dLoaUJaPwgD5pd3
qe/NZo1WPflNCYJMpqUt5ciTWDYAtUONLNQNxOZadt8LcXwlkIVHLTgU668EXQvj3fG5P4lXKrGn
/157fGAonEROTPfiCguaKo611krcKcjMK661FyDA4LjcPCklChFK0ABvnJwwLrC2leYXAep2zX9D
5becWBF54rgL8PffxE7BRJpT/KX2GF2qK//5ugG/Yx67pj4pnIJi+Aba4s8mqKFsUgHHb3fr0qmy
VESsNuUjRbYyInj93Q9zpYWZYl8x8h95v3OhK/3mckP+4R2df97j9VTzkYruS4NEqYXgfAIh4v9K
rrnX016ebHu+B8R4fvGRYvsBF1EIIinnGDtzQTNkF1benFbFqOSy8djH6kEla3s3j85AklPfcfDE
FyieVc0E78X8waN05co7wNZ+riidUF0/Oo3gJ8NivVog5YcMJxmXfOUksY3lWWe+AKOcYnrIsn8B
lHDg3aLLa2I1Fz01eLIs68gZWgVr3qHRpgFL644E5YnreqN7EPIjNaSjkhamKH5fop7VXctyXBXV
gXNaoAaRj6A0mzggUZHqcAN0xabHqg1z4s+2g3VUh6S/RYhHg58BLwXtH/icRFB2THIa9wlvYTST
K28thbZ6my6yT4WPP0Isz37v5qNJkh6/fIIOLotvnMpHDvfOzVTjzWW2Yw/a9btgzoDAQG6/Pelb
2M710I9isQ5ARNuPM6fW/+CeG+kU0gYvsyufu0D1qpQKhNqRJNDc1mlKF+QIi7qmgHlT/qhBt9hW
3v7cbzP5UhlxvhOsjzzhwBhwoNSSejUQJoJDi1JRxGJ4aB7ZNNKOB5jH0mMFY0McKPHn8+JlzkfS
XjZN18GPrKILbSF64jdDJXQhFtbaVtHtlORNbncsArE27+m7W7h8eGGWWvkQCL4t23yc4GPLGznC
y2HKPditBFHNxxPUr4WuKJ0N/RJnC2tAuhRdMkwjOeG24m+aw5ino7XJ93V1OMjbL2XIc9v5n8qi
/7oJqX+eYADcsfLtSrYNMOGQ1Q+4fAjbxbFD4snsr7vAzcAf1JTz77HSC/B+aX2alj+goL95arNs
9bthd/VMWXPqYcBLk89fV4I5TVb/7AKB7M2A/F2b4UsLnumIZthPnTKo+QVeN7FXVeb8KTtuP8+C
B0OtIE8xAdq5kUr+MXgw4Z3E1QSYnHJp13ezMINliujtkwcaX5zW2UnWevKgMFbEIGct+FJf6lNN
e3Y4jo+V3m3Q3s0heucgEWwTTbownj4jyPFXqswZoT8K1JZ9KSfz8Vr6hlGwX4oUWCYhZx2J+QD+
+osZl+DJkCSRnGiJ6o1dI6zZ0S4tGSMwUDOLVYky9UCmJGHIc3DRwvGrpR4pfdDJXPlMLC3b0N3Q
mTFgInfFEKbAX1cC792yKwlhB+Z4p1djI7es39uHROhKDtvWjls1QktXAluYTn8jD74LOzVhp801
g+WGdaxwNYvi/y58Q9D3lgL1iQChz00nrCbYL5OJOguY5RItdTwHyhHx1MFBsdIWxztws1IOA2AZ
AaPVbCq5hcQffOQkje/E17JhZ/zkSYSGxZ7f5jTacfk0snOb2qm/PBMIJeGS8Pe7uAmxQwJDqQhM
2wRgr/B5LXNc8KuFEgUSVo+/GAFZE2EJHvdfd/wfoOo1zAn9wX6+3mauF1l3O0e53zmCfNWNNqJQ
MBqi4pdBojVSKa4Eh58UmzZeG6rOERDZvRVKUGqK+kdfGnP4rSG5HnxTrsUj/+lb1lQOAYMV+RPz
Q4KFdH2qYugkWyA2/fRnPidouzKmJI+iE5Ag76CncRFg0RWOjLyYzncSlw3iEKOjNGDQy/O/Cm0P
ck74LZUWIyrXVOwg5WYXmd8levH9Fj6NfUCZf7Fs9PdDSj07ibN2engpspQXbEdR0RPMmz+qqrfh
rCrgIHq+MokcJZPhuU06KBiQuW5HJAPduxOAOXD4NL07KBxu5Y6otlnkj1EUxkq/XkC4dv1kscha
G3QrEGYzyZyQOCxOjG9Wa4hsgfO+qMzCwFQx9BesnsESnz74NuURncYGSpUXs9eNx4oR0QMYE6z8
M/tXfrA5MD/uX8v6gNYYG40ckm3nMKh4t6r267gxi8bdnU41+UjviV69BuYnTllNmZGDgeeUfd2y
iXYPA1qAsMvVM4fD3jNVrjzFQ8p3+UspmqMHRpUsyOi7eTNRNIAXwAj07zDzZ1NyEKAeKe/49k0Y
p8e1v4Wg/qfarC+lHVjbpOeK3C5n7PtCH5fXK6OInH6AqTtDpRzqRUKXIUpVVrZuvCwIZ3LWLfPj
DkYlrewm5kY4w2XnR9zdlLsxw2H39VZwifaukKAzT2WkgogTz8UsZGQVukp9K8MVv9D8GAdpfo/B
NrZKBqVyvprEyyxYa9+tKcH8aKmkb5Dkgg9YzzBlns3zpGfnzToAXQGl6jIaWs2gOzYnX9ROyiGw
Tkmjp0OGSds8t5APcj1tkanKl4xLj4yZZf7fn7fEIoqpIdvT4AHoGHJmM8AX517ATZuyu7IGtZkL
pdcs1dKqWGJ7eoKbiQST+Z7PgDs9lxeTpBoVUr7aLgkqYvNKHnOmlw2unMdgyQuyJatrNQfiJ89P
KXoXoo1g23ouncf1T9KJpxy7JgUSW2+1zevecgUKIxPPzkgnMPugBCEaP84R/6vdH+AiL6DEGQB1
B6jdVyruBZpvVB3eNOoc0tiunuUOTeAi2pA56D7W2Dtdv6mZfItYRjLV0dr9W6meouq7+nrHpfQH
admj8yAugI20CTMVanYqAxqBUE6Qlaxc8JJqPAMLVcLsEsZPJJrw2oe8s0j/fDkQ//iY91ImzhCq
xX1w2e9pZFUe9E0xRct8ktHT76PdxN661IlqfGcjwcJnqOYM86zI4OoD20kPw5Mg+dXvpiaABWzP
zYqVemQqd2quv1tRvkaqxMVYKssGMMLrbGcj3Z8p1tw4Se7YTWKw7E3AeyT4Li80TF4gGNesjkiw
l8LjzcrWNvcAdr8lAaZHrOm0yITV2437Pjh8r3C9L777LGyBIRXgi+3oxZ7yH1v93bCogKcXWNTZ
7QE7aSVfb9xNvZXkXi4Z9n/21MYqRyaRnZgdTx0LCWhrwDnRzQdZEpXRWqrzkHNab8nDVAjHG5pZ
sHpKahYC3SQ0X81/eOBABvGpnlKyS4pozGSUsY/VcwJYJXwyvlOETh/1QPUzd1SGEmEIYgLErACF
oniBNB8Z+LBRkZaiEu7KN1spvRqM1cmV6BtYEPQ+P7Esz6twgVA0xaqGwApOgZx6hxiN3i32gYIo
E/wZsCQITjYYnX8s3GvYeVQiRmIYTaxRAOXzDyhCjpcRT8/oSSY+uPh7HBSFwJtU75/vg8wI+UBo
NWN68rrEdmOwDwGeMh5jujXFFpYdMcjm+3fpe5j2k+bOQV1pkammsHRVJ2B6cY1ImDv1ayPH7C3U
14idPsmG9w66KeACIJbi5D1blykZ4NOhGpZQBLyWLdzi/H58qu95LjuNmlYOLa+TJFoDu+FnQTYV
Ayep4a9v6IpX3FKBId62ziHrW1+y+K/FCOblTys2cF/950sb1hFuDkPfo2jEvPgmT5g82/zWpNp0
5fX4+bynevFBzTHlH8Bqv9WbbiSdC021zNvloFYXJXAsqHhYVKPf9j3ZTioX8mOp58QVWGrhOPwi
TiXMNCIGHK6GPfrmbHwKz750hzTjn0Aw+vVE27F8gO1z36x9xPczFo57pB8uqCARUpPJP4QMvLtO
1NhlOd6xmEQ4l1atU9nCrJjKURdVPeCmDTVchunVOQkqYW1kJFyJexbk/QkPF1oHiXzOLo5z96R4
l+GADRY8sOUyAtHytDP4srWhkxowZ6WyfEoGVYwAOfIxCkNLeNKws1CfPNyfeoftKgwHgaor2m+6
RbwXrlBUGys27CAubo8NCpU3TaDoQchqFvd4H1GkTb4YLFPfNCVAO+94LlxtgNBsu5PLyuvN0vcI
GWp16xTEBaT6/SNUrKtB8KkhpavG7+xwMCOIWurJEBnW36fqQDgO9Q4vykfJTsIC6H0dG2oK6KGH
gowhcfHOSDBMOVfq7at8a2Yo0DJyErbmlfiOY2U7Sha0SFrlk1XYSjgQPBHMVmrepmZXo1jSwm99
EuLaC5Tk3CwxE/jkb8pAFHqBlSeT3Ake177O7InrgkMT5yuzP9D8XhO3FWwLjOspDgAIIDheh9GF
sei9e2pBqszjHNkCnodGL4KKqLkDRSphjOPosWwlfr0v0a2MhkBjhVuJNDqoChLYP8wPb8lOMIxk
zFGe562QFw2D9dD+EnklNpo5RQvF56UkRk8oPlsH6jYpkEweKbptnsHcSf2fsLgHhsATFmYC70B6
Ro/kOxbReoSXXrO+dHdez/P0qnNNKbju8FwAmXiIrknzjj/BdKfCLTKrxMEc25986GAs0dhZnS2W
ubNmtD7vpFcCtB/m6WxUJ9VT9w236e7LqrBwa/yoRnDoLwxU+pYB+RNGM7OW4pX00vutybncQW5D
8aPW7MRh/tgHOesJ7zeyXRt/jaQMrHf8ccX5htrnw+w+0KoS6g6iZA3enIbBbklmeKptawFKkpbm
+upyzCbnjymEhHQsj2bmNrDel9AUNOUcf/twkUTSXHNyXIg05vbyKkYQ4Oj2yl4Ev37O2hfcalPC
9q1tHu5Lb4hiz/uQea2iLinA5Xjx5I4MLuu9O8gOBM+ETqDAkILPeTrCvpPtCHMPugd6SyvS4Ae2
65v66DOyAl2ssoavIUopiKpvMCs46reSIPb/BTBNrDl9Fxdu9IYmsZcrD+uRx6xC6fQgWzw6ixws
K1NNUf5WjKqeWApik+QagdZBcPnfBIVMWcNPwtuMmP8oafB73U0YHGh9D45rue2W3omNftbO4s8u
awiG4rl86ed3FT5jBSzUjhYlCSpSogjzV+fLWDAa1CxZioCg6OXqE0li9mWZ6vgn5apbhtar1VKz
S9P7DG4LtoqWsQqV2MTKQUzfbDUwdoMdgzWIGi0AUI0cCZqja+4hoRJxSKaiQm4e6oMuH0CiaFgE
CDod6GsoH64o9eTLcoO3rDyqvrd42JTz8kRuDdoQgYziFMtD5MUtnmLxzc4PfDSgeqpxhe7lGDH8
RsTJS/33j7+6sa0f9r2YPTsT2LGPy5DGSIg0TtKhu8I7lZ8L80roErQ2G0tfFzGYnmT0QVRug2qE
5c0uT/WgER98huy5+BIcKtnZxzDieJ1vI7nXJvvs0YaAu8KsHDvUBzp/kzQ/BfJuUiWqkkvEiOCU
etBHjhEhwfl2wirttZoVYQZYkeonDeb4/VzoictD8gIAmdVohELOdALZkbM6LdDm9llxhSu1+lhV
h1FI8uEgbDRwE8LTYAqGC5V2uQqJsJKTf/p/r1ckPsodAE/uiLDsSraq+NQYEbjg5YN6CsqTw/7v
psg9IMOiCSnu75JVigUy+lS3i8o4C47u6n76vkAzQmvwCDDEmGz2i1apnn+ng2WEO3u+qR90Vnpu
dLZu6XVe/A1mE/dyW4tQJ+MPb1s3dWTXoLXnjCiTgUolayEBz455LQQMS7NnozPy+l8oMw0detaj
snsUzyMQkNYg/bXKOW51mch0zcBertGJ/VVGKCmYFj4lqkjBB8EhqVcLeO4SG+nKHcmj/yw/ZNVO
FLSJzlqOGR12sNIU+Rw24iJY7kS6HHWTOFmq0O3orZPryQXoYD2J7NnxG5iRDOSBXBG95Vluuvyd
TZygPSzX/7syrToPR4f0SYIhAaP3/XdpGxM/Xqsgw2FZBkVe2ivExFnHJ3YkGZqPm2/flD3W6qG4
DejcMlUkHhQUJyJ3fe3P8NRZ0EkLG+FwcLKe14CmTtghjnqQhRkK1ZfXrEZRfHRrOHwe1Z1GTXtV
5wEGgynbqFdyRh/TwKgE6YdHZqxEUueIBBaqd6oVAGtN29v8UcVsdt2LaooN9wzYD4X+Q35IfBBI
Sj8QZoZhPFA9oOi31Xhv8v9iv05CN/+o2sjNQ0QLgG3gbUISAMm42JGZ1MOt93pDUlgBGV5RFCJs
Z2jVb9MptWMnowW/OTkkSRxi0FKsqUPGM8IZKiGiAd1MhxyJkG9f5+Wj9Icy2onH4LWNq0Cw+Hgl
DZEzb4/95LAwzZ/vqudsJB6EslR+YsaM48FjD+MRssGoI1dGR6Bvq42Ix0nBG2vCqA8KfuoN8Dno
CBw+fX6KE5LP9w5cxFtJGPLCa1Ih31F6ZqCOUdzAA9Avmjha2SoBFfq6WoswuQUr+snkMG2AeeDz
G95vsQMqJxUUkvEytaYJLEwBpEOGEUwH2tv9WST0QoUyPqW0yft1Qsju1EWEEspgH4v/wQAiiHwZ
68r0Z++NhIz7tFaixD2LC4UGFxzuJaf9Okzw9dBTsEVrLcwT8nXzVup3avSJG6aiC2ssjmM6GZhe
PHHpAYmBgglTyHZqLCgnh23X81RfbATfaSMbILloNb+GWUKIkBPzj3aQe3zUm2UrzjvUw3JtR+WV
A228P8snIvFQt4KRWkJjqejG3puxuSK4yWeSM311NyTqJYclAwHwTIILnqsl+xIsZFrduWZJjyQH
+oO//6utyFj993sqqr1WPl5dPG5ga4o9naMkwwVOOUHQzHaKsQu0kaH4czEPiPn51Zy4EJ8MklqM
Q/R11D0Boe/m4f/wmr+2QB40GuuXv8zCB/lo1fUkzCccBRk1SVvsFrz9as3zKu0j64qIkrliJuVu
VvgfOFqa1+UgUruTg8/x5dz55pzvgrzwvfdgcS0vL71ReFcQrtjs+TUxlPKSBNvTpfgQ1xaEuNyt
G6uRUC1ejQ6/WC3gYIH3ycc4jp373O+YqW0NbRLzvctgigi0+M9vb/sMcZwMioCiDQMGaK3QkDmn
7FolLklb/ecwztE66j/2TpXmWLlhWmk22h0VuAanL+nwj9QqTvjaqD1Q/qsVBSj/hG5sdodqwKaI
kH0C/Gm38z++dIq5Ru5yIQYni7M4gbnvG9zioX2ASmIlCpzbwiP5ntdmzumCvdVWtVCYYvxkvGBU
FyeS1SrnbuEUlP2AVwOzpLXNO3RBuzCJ5zlwjp+p0kgmR7D7Jxdeeha5bSid+YGCmcp9+9X+F2QR
eZZ5PNaTtwtLP31DWSbu7Stl/iqunb4cv8JhBQwTDxSehsl1wuoWACOj7RvKn5/0Ljx8G9n8tQ7v
noia96M1jJy/6FoYiOiEVYZc5Hz9I/zsI/N19Ov5sXuaxYAZkW8qVPafoQPenPEUNveGNbIyKOh4
vyD/Ij7w89fPIx5fsb7pZq/Aq/VmrX2JyPltdvJsVk3OqTJiJVlCXaptKJnsEGKn4b5BPDT5tdog
aCCT3DP8ZTuhda9TwpjmCgDfSmTaysDX7jq7EUQ+jQXa26pb88FVTFt3h1xQdp3s/pWIWNlnZFuu
AlXKLvAKbpyQlBAiBZQuiq7odLFMnFCzz8l26Bx9+/U3yQp1pME39aAo7/p4Y0Xld1F88EWsVAgx
X5t0XD0wTQpAlJAs5eXU3ui0Iw8htPwuX0qYlir+faa8lMYm/qLLqrbPuRbnQmyLRJG97zChZv3T
zlFKMX2dmgl8A4PFnWoYJdfuqkPnOIepPTSrkc1WKaEvIxtLsDFy7MEqy4rD5qa4EWgJoEBU9ww6
UZ3snoWnlvIs2u//eJpuRNeEiCw0LfDwTReFty9lNzbGPIQJ1v+3RyUrBZwQJuJuo/VoKEcVrjNI
DLpdi9i4O1TaKskBiCi9XZ//TxanYJ8l1S5W8kanCqnyZA/lbVca4htPWC7jcPAiK2r+/dV0rkXH
SFLEiB48PFbHD6QFeyBgg/zgFohSxCr6DoMeR/urpx822Xu8ZrdRYhndBIzBf+MA6EEeuWXTXHK4
b397cAWUz1mjEgswj5N6KGLougvVdNqKSERnq3X7OLDfr0iU8z+mixtBy17zjcArnliCJfYrfZQY
9EKaVTXAQXkpDrfLYTMsHHZ1tM9ozrmgZB/vb1sxS6gHZi/Bq+rk4AMwuNi21trZg1W2JEq4FNxz
L+PKTSCp2KHspHz+UGfSikiywABWdicZcB5tQ/XwHShr0KRez9CHHdEyhImLyuo3N7km/3paRaU2
QyLhPSW/UQwDs4Z4VSg8rcK3jDMJ1ydSCrkrhmHGn0K1tlYoaIb+4faA1aZhhIcbCS68hha7iY7H
+v1gnwwIZSYdtAX3TNFOOu3XUKBC3627SZXOrTeB80RLsti5ise9dqcL+mzAOGWnCggzzCrrWNZH
QF1WB8pWjcMqh71FXhHZP+zBWRlEfftFwS0Fnp+w4lgNnPl1forhEqMh9X5Afj2pTLUTFdMNz2ZP
C5cSmARw6qidxSnmkR4XFXcFsKJc6cXE/dwY3Ax7lW8PepumFTP1vPPwHHZd04uXm1kSmduwszA6
udsNNQ1HdiWgYmk9iISyaFIH8kCm4hyrVEJbjQO3S5/sVLDrAwX2nM+JLcKc4ZUivorgd3Rz3Yuk
Xl6Jqyu530Kb6rVRHGHo6caeHkVWfPJjBtqhFWREm7YaFscWlhS+/hN0sucb+3W4p3+VhFN914oX
s/SaqM/or5orGeaZTIcQXh1ekZIN9T83QBDxTPtjI0IA55E0cg49ht60yn+F5I+iRvmQrgYTEskr
bHr1biuH6w1XgSGd+7EIuP+pZ+Wipt7glORWN72UnJFmYDYSicq2q1mrOp7mFL71Ox3R2MSA5oBl
PwMY/y4h82S0/ZLJ5or1X2pBFWogCc/3vF2oBqufp/vUfCmDdG0QXX8wLyL+boTsrVCnwx+NSd1m
YcjzsCr5odLtSjeDTGfp44sK1q5Z2BLz0xbZCF/HkraQHrGEfGGgJXAHsNOncncmlLWI/UkV3J+f
LCBtM0p3nYqNW90qaNsOdX0Lzialfq6lRFitS7TR2WrVbfPXVuI6Z+QBU1s284J93REoQlY0btxr
4R9BUienn9xYdVsrFB4nX/7qWiYmW4LLHX331vPr44hwAetp+DsgGGL9rI1zBH8dXrNWSQkTUCb4
0sDzeDnnx61t9CXsBzc+LrUC+Yio2BsvFDYe+DHE+n4yzEr1GuvilJzq6+87QYH5lvqbTQ5Nb0KH
rcZQhWcKLki53haM3KgHrTmmj74iutGagV04f4o3o408m4Jvzk6duzm6rL3VM6/+K4ZnmcW4rld7
5zHe45wNfveHaMywCjoaiySeC1sJeLauD5+DBx0DS9xtkBzH1WGUZGo0U7j8rhBnnWO4QmgW+fvT
WzqmxX8U4BOTcT3mbfmPhlnBfwUg8O2gpVQJTkDkCOt9M//JfI3umPgH6392Fc+jbPaKwhzjb20f
GS8SeeD+JQ/W4Zm9NmybAsiPtDRdVyjDRddAavQNRhhYHuzlY/hVilu6jeJAHDSmNwsVlRgDhiMk
HiKaWgu4oghYR/hoIvQxSdimpWSWCV9d4uB8EcBR+g3f+UU4lofTzpELRV6gzav3h+2s1elM1hTL
am+WpygFnk3peZAKecRKnRFJU3xKNUEc1xVaJuN6387KBLX/t43YX/BUXxnxtlB4pc51PdnwEJLN
y56cJf1aNRXLsrcbQHYfTzRHl2c/XR5OP7q5xp6yh8Lcc/7i9C+N8h84IiohgOS95lZKPl4K8Oa9
rMqrC4uW2X/E8kDDJ/Fcs7DxEZ2vLZw/QtM989TCSHSUp77h7G+MjBlgmNkA+ql5AjksuEKRUVGU
M9/3JGLzdVvRPDf0BFyQtpnaSIhYO2af0kmwiy6FBHAEvPUw7+lNLcVfHBb2jA7sAKC51PAy4t/g
xPYUzbeK7qOBP2WlrWMHnOjmuf0x9iLEZ6qGJWpWAY+cTlnUDBiSYAL1ONocjMt4gykhnM6bjaW1
hTPDcliFjfs7u8D244K8imSh/CPZ7zFQolfqRhjU8BntqvR9mzF0UQL/elwlu4dtTqrGQJRo53/Q
hhtMSAj2X1uGxtziHx26lHEI1RbBwwc1ZlO/kITEDHdfQmj+pcJUH2oW3M8/dzqmmIfoex4y37E4
/bdyIKhdskTmlp8tnjLxmsyNlVtC8rg3BGqzbgK6h0WLhVMFOaw8gpI2S5GsV1qEce0WhvaSqRwx
J70YucZhDqiO1ExlHr9q49VXvogl8rl2AnJvut2LaeEj2J1vefXbYuQNju3Q9bTxhm+oc9rLr4Kq
YJj8z42FSKe3K5ME3woF/3lSONPuY0xOiZFFS39vo6Zs3eYw/6AtOFyPLV651UOaONdlEg8AeP0R
AqQgdthz1FBV6ChtyD0xD90ZtEpIlHzsJ7eTCXalInZsi8L/gNV9CUzQcex5XaIUImirUVVlCoeh
v6dycYRs16eRMAP6YadStquOovdtJ460wxz8KE1HKa8/mxy1vTBmWon/kbwjmPum+3q9nV3u0uOe
YuZkj5x6KZqxFWLvmbTHBuHMtye84QAYjMQuNR/9kYVyO4YIy1wifgdNnbTDPNocJV0D/s0kiJ9U
Qzc7w9CsPcTW/HPBpXTJND2wSJb1IYZzCBdeln9+xcrgGdptWbu3tsOHgwSN1bRz0kAcbRIwo0Vy
mT6+GIYeB6o8j3AqPUaplohrDfv8+ZJc4BsROKro+VlZD0CycOxQaGPiwDXVpTtLHA9e7dx12GxQ
U+XeUSNTxC3+uPcXKR0X1PIy110gH9aoxe1srdVcmPWOE320HO7eJKk+fVdpGRt0o/STwgI43W0p
UYXgZmL+C9kYMsF0wRB4M0X1lhCPZb6JrCpMw9TUCKt4QHZCFQNZS8Q1sgMz73OWhXLoHpZwhrGw
kM7GUqiGB69hLWPVFcXVn2PWtQjhxQxOCUXFXL5ZhFTzyol+NQQ78VDjewnbt3nj6GIMQT0nx5ib
BYbXql08ea5QLFfwR3vE22FUEJlJ7avPAPlt4QQ6gILyrUjqQq+NSWtN6eWD1rWODy7LaB7jGT/D
dThlyuZa74jUsh9qKwxYJDOqAoiqfjYxV0hBGCpIAq58APl6T6ys1d7OVezcB0Wvz/eBkRYqb8ZC
tY5Ze9vPHFAZ6jaiSEcgkj1Knuq3aAybdruX5cpVkXhc0bedMFWl8LKIXb2HwOBpJhTM6z3PMpbi
Pd/WSrKL8ue02fpsnlTtHdqyo6IBfNCdF4YfbFsggZ/oz+V/EUW9Dr5LBoSFUrNj2Pfk1goj7Jme
ozqcu41VrLzbPAAEhOxOIXMPYg/DYtnJCxEUTe8UD8jAZfDqx5XzZElYDdBlkSv9eEfGrl6X76qy
2NPg3v8WwkOmEyoilBRBqbX7lACb89JjiJBFZIh89HWIbqXXlpj6HPVZesxHbInkzXVFPmogVUu0
yW1IwdU51U9iwo/PH1l3Uk31BXhUGjFfO34GBAYLJxJNI1p1c5ckZ1d1pjYod7voFOCCKTVYE85e
BUzg6Jc15uuGTSW00iEhHCiCcAjMO73rK/Iecndk54MslbeMEMGwnN1F+QcfyhYHI21wGXpvF1hE
i/8k1fptLaT5iAYxWKuK0qSuuwh9JP0QpGGuUuuxJVqZBEqoFEamNp7jstlK0DqV65jS7YTg/eTS
yMSGme6bQ4dZEGMTWa4RiBvzHUyps//hYoo9mNUit78dwFmwy2eRtU2B0k+8FJFR/wlW9F3iV0UJ
0RafQ63uKifkfMDlMgBz7ylKTd167hnzLX5CBmUSEZTBn90emnG8uuqBH/AO286vMsPyhd9E29TZ
W1FXO7pKtE3CmaMndQBf/PTvKKFIwuNB75/pqTVAy4Dkv8TVK78W4D3KyFmEvvISMul0qHIFCScY
2/i8RhVUZ8+Vy3UqvxNyKqEBO9d0tGIbst8YAy3gVt/haxXez8CjRZxmREjT1dFmZIQS/b5ZTHil
0e/A4Q1ccCqx6aNizo9zhEnvfwXqi/jDa/0Uv49mUw/JfyhlN7AuWyv8LO441KHT1L8yJPPNXnMp
NDmzgwhZnm7rFcAg26Z+RJiN+OfX2MjfJ+jVQsHH+rLLZWEkigZq3rL36zOhjgVgrwULTUaDgMWI
h0w/Iu94Lc02d1OlZ2NV7cjSzAA8OAhdUfJYfNdIcBv467yAn4XL0VCGxWxUTB4lo+AF5R5kn8m5
zYOTkR7y9jRCmFhILXnJIvN8Nrf4QIkVZP91KL50UOUL8MqNDfDQLVzrnLx6XZ4P7+EYt5JdOPG1
ESqTMq79gsdQpg2ntoWs4GOGCj/TowwExxlB3HqenGBP1fnjal107PTfIeUnrWdXYW/IJdaAQxZp
V1b3Erz2peZAHcK1i+rroZiFnrK32VYO616nyguidTAfa/F9/zxvf2hhSRnVKzc5WwPev4ze5D3X
NF5ABXbTnWPvBqwYaI6vmH7K1DKt614LM2V04FCW4yTn+QQMDyK4uLz5znkgO4W6+nuNoRcluaa/
9yZ5bpezIirwGmMYEtsprFE+U7x7shzo+SDuFiObVRjlYoZZFEVhZxRWGJJSZLl3377bdCg6+Oxs
ueKJulAhWpXxIrLfIqFnedGfO0MIv9MH7Cq0jPMPeZ+lX3yeKHxQHCnwOe31v0M4aAskUVmheAfA
DvMPM+yAnCO3nswjFRzR73izbMfJaVjJ85mFXyzBKfMQRpvVeLV3VhOY2DN3Y9eAhTD2O6a952Le
nl/lk2f3V0c7qYriLdn51pzYbNHCPfuz65ACyBFst6fdov70d3QxG/aH66eHxH7S8XfYKN2Lkt3g
/zneOfkUc9EEjN+oZcEB5J7xYjVHkKvWO/cew+ytvLbyBvlzICtlzoVyX+TVS0ywDgqnv+ovzWH8
IvPPvqHh7eovz9sjaLN94iQCEbBHpfIxhVU3yL9q1q6L6gDkl86+KcrOrI+xKSWTUd0gMS8ddyl9
3DPLcoaKgLbB+16KnbPi2BWOYxapP0i2E92aIbIsc3bRtkY6Q8i/VQm4h+hRQQJLKgPW4uPqSov7
yrDjOxNXmaIcCJg8tenLHUbaOUFhIBncuqzulz2XH16ebzv3+nTLEFuZnvCItfTg9CfoGR5koxBV
M5Acj6cU8mOkZYUVkqKr4yb+3zNY1k1hL75VCFcsiLC82v4GgD/Ji4gmiGasKNNQE6uLoP1TpAEZ
eIqUtatX3W7I8xTAh/ek6eOlkaHcLU056LWelAPzi06tNAt6onwGIn/vFfmEz98S9bj/SXHZsjPE
3rGX9viXHs7iBW9/eH4pg70t+a0fKlMgQv/u1Co+FOOVlnnNxnO3qm796c6a8zWY6nED4Lrg9AL9
BLFuWmk3QV4ND5yVvAZGHHEtqmgUO8K5onJmy/2QBx6u+U/70dy7F+lGkcEzGvb5wcWMNYu9cxXy
EfVL3wDGldO3K5DS6mQqP/4IdEjUeGZs1uErIPECjeuOj6sp5Gy8uajTqv2EJyv9TqIMEt4qE1Cj
mur4tS+vCdhei2bSCyQOo/+VTETngvDhefliQAn3qjwUoQQYDs3eX3cfUzRrYIblO8oRFI3RhKTS
b6efj5kdv6lNBbt1Zt4AmKwLXwI8bSSWmZgZfww0G4CmyAfxKqDTuMWmulzdXCKBHf3wxSpv5ld0
sDTYJgWhirOZUq/hSP/6ScTfG5Kcc3yw3igiXjh5NGdQ7sGP0lXnX1bmTvaGj7YHiSR9756PBNdX
5HnWMcpD2AylOoc2jZX82KAnMjU7NdUKbuwjHminwxOS6KVmOmJacPllyuvkXFrd2l8awbAGrHXM
18MMvzmkbDBUFjhRSjFQJo/020owxBu7HqdFwIB1QQn9BiWm3OiuWCPUhoPPs4aM5gUNczE3V4DS
rT7RQF96FnRexpgdeUSW4/hOTs/DrgX+DwHX7/gk4rPhNhbt2wFhYrplsn6JnR2TfcvBS5v5CHgF
CEGwYgzqErUdluvyhW7SsoErTmfSlXioIX4GNmvtuTMcBUHZ1uG2CWV/VSw1o5fPohWUXjjBPw6W
tjHndLRDm6a/HDXuWy4GEcvasQMUfNbIJ6dpA/hneQH1aiXQbko3g2/pquZ4SaJATgA12W2GETpl
4wkjPKUlDd7lJDwqL1SE6gn2nIDPTdxqIVsGCRvWNcw8rEXs2LD6qpPagBTd4yLVBNBaOqYnTmP5
xbPZKFBoi44erW0EY+iVr25FJ/ar0/TNfZRWG7YO36uLHnvqQBrBcMy+62xkD2OtBCGCZo9ADTNw
gczMTvx37qiPnW2ZnuRbblOZDtVQQFREfzojn00ZEPOkkZAP+DdWkX3DtVXoKdf8EoV9L//DHV2i
RfDO8fLPxce9MjtcfwjqhfRlZwiHiF9uWl6TaUfLmfuLf5PWFkfdm0tvjifgD5tf+TfLcVa7oThv
77UpBqZf1K1VxKe2tkDS4bAm6LGEdIQcmSypEs5tPI1sd8LC9aZ2a5ZElNwlyEJY0+m10sihsZwc
D0rLz/mwKIHedXi5aNtccZE5AntbFLYqPyqxQT91TpkYiusAyhqXfLAJl/t48XYUR/bZIK4aXacM
8mXWDsTscxDiQBNhm0ao5X0VM49yCDMYk3ggKYjTLNW/LkZ1RX0/bA/LDmKpCxcSEFC8IK2HKUId
OYnXy5c6S1y1Jq0oi0MNCN4g81y9YljGacAUJ6d5gNEjnf2d1LSiWBm88/AoFZV68YFUDM5O5tSA
ofuvsY8vgsTVjvmfCpcUx8/UUlUU6d42+T7QOFEHd5JZTJckQk85KJAGWvvj4EPnMTzffLOFO2i2
1ztWz7S8T8o3mSY2GlEv1zRXU6d5N8Mc6V0q4nl1TmnI8L5fCz2i/0QHdyBeIkLbYCRYGyubYmke
GeSQqTqdzFlEcimhjJDQ7HCSgtWi5LF2UfNxUSxSBPTZW2sMU1juAiaVEFcupnwi3siGDnv2eYqS
OLMlheodBm49yoGrxXDpF1bhuoEd7QfFTRZIgN/UxZW1nwEErW31BnDqBGKTJ1Uk3e17sC5bMyKN
4N+HV+vEnUqY8TcoByLBs59uGXpkzFp+eKjpaJ6PuS9YgdasaFwUFi1G9zLuc66995TfNN3PtoB0
eb5vGVwdSv0LvfW1TYOdVPW4Biapb/jqWvJ4jy6hkat7Sa89lzCu9dj0HuD7H/xk0jX50aVycwYM
kqQQunUX5IghZ29YrFgG31kvRWFgL3NgcpVMOV1aPoohFUy1hE/ZJm4G1+TZZpKkoPH30/kSqLSP
SHxBaD5FajpoZSM2BroznU12pD+jgibwvKo5wyWmk68hRa3+CxB65VB/M6HbS0bfsji9HIAm1S6O
RwszrIgPBw/0rZmpc4nMO8tWLd0euCN1UPKEOyEZ7RMXsP8ovrR4PqietQNrdNLd/ZxfHsQxZyGK
yYMGOymzsn+i+gmN/urqO/9T/MKglIQI9+7mtu4v+B5+6yiF9Kx+TngBwNn24+X/vrc6WllfHpVF
Y4PVkWggP8JBAN0vqNPcD5YTQ6m/xb0H4CqWWWjFT/U3HMA+46MpWY2cjbWM0zd/rHhlmfuvrgPs
p9FRXpyaBmAeYDECTXlRbVhMXRX10/KOTmcWpyUJkD/6rq9S8e/l5eEZiGCFBntUHzim+ChSaWxT
cAAqapFiN0BjeJyajn95EwkhdY8TxQvHlZyf0SqahmpS+IYffhnqgCj7J6/bdeosNUyG0dvEeBEH
WR1haWKLUnopsPo2OFIFGk7NgdWatp4xaR/Cmt1NO6y13sPjM52o8/7HM5gORBByUWcrNY+0/06A
AV9epdY+DNe1l+OCkwvxPRvBHmajY1w6ZC93LyMJwlLCbQwT+xB3YRCTdtAJpsi1GPiokwluWVhq
vgnG90lFHq9T2Mr2JpF4/2EyfTRiuPsXceO55OSxsH7yQE5YAIzsm8r0eH/liIjK7qx/K+7j8bmX
w3QrTed/n3ReMb5c6Jb78yfKtuZMAk/lwsjYBXBooaBoio2yUD1sTVf0JWe3frBVGJAyUfWfGzd8
xMYMcmGtcM9GPSC81QR9rLw+4waidjn52QPDqupShjKnd/emx2RyfpDxD61OtTlu4E8a74elUs+S
IVxFkhKf30RK4yg5WhNQ/Y9Lgku2SnYXD4HYTNezFa2yged6ik/b30HBQOlAyMORIZaxop13xaA6
zxARUX2YcgE3Fml/UyJRUbqPvTiHx6nj+QlSggyXRGy+IsYUL5GSwRn7aiX9sTc6yrE/7yaAEcWI
Kp1WWBdaae4yifg0uaPmQkQpF0q19v43ja79TBeAUyQzk6hafcuL5Ab+x9u+11HhWV2JDnKt82Nl
qwspZAyb5B1hB1N/p9MI/LqCoN3QHVzNIskFMKQlXKy51Zk6u5l3d/ecRewoYyDyx5ZwpOraX1Qe
Z8bmPGrjMNnn/Xp4C6JpdQcjAxJwvclP2P/fogM8dd+totFaz5QxVaCLHZLaqNVYOTjHBvBD2gs7
Pu8SE4QhxpdZFxyu6AKStEG4m4dB/8FCVwiDvQC9vYnMqcbWoKvwVJvx4ioukJH7U2/AuD5pAEMk
T29iG1qa/iNyinD1BVbNO/VuGMmdF0IL7/VfVDbUVibqzcV58mOLXsCay54HQgeXAeD5fTTucUb6
ePS1hWGTv23k442/JffXjQo0W+7VAF5UGvf5tbhFRY28f2PWnBH6aOZAUvOgcFN5GrLKY1ekYyUc
JZMq0XvGrOqYzWEwvljqHDv8Q0SC/d3NlDjodhTzza4xBE14JtCQoBGxzhx+slvVN2+jUNpzZ4s3
T074cj80KFFu3YbJHLxX2rPoiswGo2kel9788DTATP0tuAS+pKikpY6a+Q5INLiDC7X2yFKPWd6X
jxTRHXuwhJW/rgRzi/Kztj1n1WUvFyT9mbgfxSjKVjsxxnHAFGt3fBHKQMun9sWrFAgZe9aYEDsJ
4/6pwLPMTfDkY1ew4PkF2IOiQaDOvM4aApEvvwGR4+Sj1PD4vMwn8oOkTQkXxz6bKyyWktMnTNuJ
w60o3RDkrMvOIh7zPnHsQ9HloaTrNkInMgBs4X8rwOkUxnZ507HQpxe+JB5qcyGjKYsUIE9hcHpI
tCbialNXNu9idi+SGIXYGldTDpvsV/wdGrs+c6Z7AmtmiLg4iI58fKF/vekeuSEqYRwIMZNyx7C/
VWiKHhEytQStseK/W0yO4O44D8HQbLsDmulK4NoaEiLSOK6hP1eoyDn6G0vS9PdMdRBoCJZXHcy7
qbPjMbq7yIhk49CsapXFHcqwUwg9EPRzzkq1nxIOSznBCzr+d9h1xGbikSO84cKMCoOTADL318aA
r74JDWgysCk+5DcfNc2mhkqYBSr/OczIzuIwvk8JBhSjb/6c9NCI+z+/8Z2u1gN3AAWILWYWDzUh
kKP21q2pse95X+ScYxf1WfVlEMgsCqVaQnzBfJ10mGBYimQje4uSrI9upRWXWxEzTsV6SzXnXXqY
qPhH7xSeMHmhHlgz3hrvbsFRcB6KHXyvhvj8vW85F3484Huw+XUE1op4EBRmqQYrHFJ/RkOr3TRe
yxToeeND2QafXB4Kf8TBbeJRCesvm3vUGTxMmToq1Q+QjiyR58uTzsC3DnW/alss73Wmr5DoABd4
9HGkKjHGFv4GokMvxPfBGU41+zixspCltC82qh6dRqrA0KRHNw/OvvmDX5xrDiZ6D4rjmvPVBnxA
tT/XVSsq5T9zXJJuS2tFUKYVrzij/W9isrJZUJ63DEbDcH80iEbsdtYVimg5+IwFrbtSI/xjk81q
XcJQtumhMs4HgxqdzBe0evLWwrQE9XVVX9BTi3RUKSHnM79wWVJ0E384etf3z+KCjtWmYEXC/MH/
KTZTvCsmltPeWsSTLocbwLJ8MSvIa5xNyzkM8u4tVK2cmUZefqqPq/Qvo2PafyuEnYp05C4uxHWB
iiVEj7Mci/crrK8rFBSvrO1j7c7m6h15y5FAFYeqiU2SQTzwKCfw91IzVgNvXYtqMDpJLmpRzeXk
EK2BweXsO2VJ0q3tWZuhN8GenCLCkOJeqTiWMv8txH/OUxjo8X0f4PYzmIV/k33ElQmUK6h7F0bG
FQZhXqxO7j4GnBi77qMld4Uqrh2LgKWUrss3j8VhylzeN6nd+rxYCir8O0PBdP6c91EENerDgmKv
GZ9yarEE81UutpX8OQJxHVk1yonF6j2Kp2mFeqjKTQc1HnU01ykpyIYxwoIifC5eZbjODq8pfIQT
SAy8ZsgNUOgk8oAHmd9p7jRhu9M1bOxc6swXwY6nX1fjGqoEqEiXtGrBnsz836bZz+/yHTAcDxJY
s17d3UPr4p8OAr0rq61P9i8WxHvOHbeaxjnftpu5rIepW0esFOVdtoQgo/88C3O/b6Y7rNPbmGzX
lmL80sBswlUheqb+w5LGkC0uj7xl8PYjzN4jeC/CV5p8PQpgAwzAc5FqlAUcPoxjUGMPf/yF6vDV
JmzC3BiEnucGfKTjhhcSBmtRkwh0nVn97ooQYvxwdlRS8MYGYuLDd2vbTNrq25CxwZZ+AaCy9bui
ig4LJq0OAxeLotbxD6rfuL2RG2Buj9DRgaZkFjSWFjgTQDRU1CYWIKK897X1OEgEMl4d0eE3XYq3
sP57/v/2+mAwmYoWHTL+lNLjwhRvl+q7WTPrY4ZT5ETgm7KiqmxVbF5MAdyo1+YdNhlS7p+HWeXu
Y2lbOSG8FyUVcRDLB4Vtj2Wnqi8iBHLVlwhnvzJtl3Y5H4tO7eeP5NguUUv843whLue8Yf/eSKRD
N2xtabeiOwHMgc1ioYQWabTWDtQ3LFI18fwWMQrBvHzrGT4DLJ0qIC8rUzFXtYdSDcVdauY8fFvX
pchimTSVpUIs8o4OtnFmAa9OCGMI5f/yz2jqHHSWJokJnXUVk5kr3ey/NoA79EFaTiSqPZAsNw7s
FROS1tMbkB4ehVzXKms9u+j9rktDkCK/0qYt4uE/u+8UQc9j/UKcvnal8MMCI9Q81tPKx6oL+/fu
sdLrmm4aRd5ekbivdF9UkP2U6cK76M4NPlxfUayOY4mDYo6Zp3Yoz4evkJMHgX8iI/CsWnTmPpUC
YvlwGPeeVaWTkOpOUj7rzEO4RXxSrCDFTvCCTrfpn3VBtVLzhzmWKCU2DdY24Up22Q3nB/eGdZcN
tC3T3BeCLiht36sBDicKWb3rB+tirtyN6pLX9vHQvy+RVd/mRgVWZYOrEEuUj7770sLn1mnJlUUi
xZFStHo27SX8CwJpqNWfXENuhRj2WjcJZMLaDdo0QtfrwFeYMLSz8hobYUH7aBVEaVsb4nCHSPYU
xFLPaxELT6+dW/vF2amQW5wOJQ+qTeDXnMf7zHriULThMH8adp76OKndgXi52O2urRPLtooTiA2M
puFCnpqJdNCghuKBqmArJPzjrHd73DHn5RjqF+u79jGjzj2+EjXqQK7kKVwUmd51kUgHsD4BOjN+
dIUhJmWeh//NbQgQSgy27pGWdv6HvYQHFswWZZfzurFqiOFGY1IRd0g8URJqfApccpwoslY2KbSM
EzndZ0WbDUr2534OkAzDFZ8ecwZb55737zdwN7Xqnxyd6xiEVzGF+TgG+tkfjDmHt/cgLSH0CRdZ
2b73fxFFw0+7JOfe/Eh/YJ4hOaG5Zu70NFxiqEwZUlptPLDnMP1s+TJOeqpuAKUNbiS5blBcIs1w
M3eP4+z4uEJ0sYid4nG45eWi4BGe4XoA7iTFDlSkyrNz5NVbbG5lTv8xYYF+ZNJTHSlEdlVRK9Yy
/Ya7ZpE04rFhVY1ebtvW1ZCNtAFWoIXt0sEI4Q59Mx7UVrtqE9QA7Zbih9UvfCyjLqRok4vHwZyx
T12s1WSZ+RftE/XTbkvo5IQVkULQTiHBoxuQVnTIbnF+wLXFsy9UU1+pEvcKawrNLO0rbJMpoDbm
+zXYPbt7LaboYWcceC4jkgFAy8m9T5X5OSpSLN6pRTtaWaC18kAoXfqLeq/4YqT8XB9sIrEVwIuT
iXCFDYpKstk/PZAv+E4aze8bwuVDWnMr9VOt7sM5YgxbzpVnY6hDmYDEWGCSax6jfq9z4t6J2xUg
SwzMmnpajdOif2jRd6CVgkvMyAHbqrXVpuqcaf9mjaXINLp7tG0v8UgKgdrxMqew6SnR00U4NqGW
kKAt8z6qAGNCayNdYzoC7P5c2O+he8Gy9j6EDqNVEH/XCl9c2223bHHRO0C9YduCWAhvf+JRfmhj
UpgZKPfKD/QDFvUZunx0z+cf6qBxsRPOTejP1JTpZ6v0/TtrKzJuG3LqLr7OVu0U9su8Vp2B4O/3
xK5PBuBP5E6dzI4MqPHpwg8MsOgTy8WzBhDY0Ff+994OoK6bZnvUmAa18q0VMZYJt846P8mEEqD3
hLU8FgGPfWUsGCVDnBd2UcR0iJEZHmLo198uSjZq0+7HI4ilaC57MfMhhlfsavfiNgyRMHIujnvx
XzC6HtkY9BZ9ywCIVl2q9asduxdUE8+i3t2AvBeMefmDmYCAUs1Yc4tTLMiCwiwIY0hb3bXjeWXa
cemIou5DUVPGFmKQYT15PO8DAfi2C4aM6fCHI35nz/WL8Nr/41j7oAe8JX1+XSKt0nJs+S+5YNqH
kABpJQi6jxrdMhQGV3r7NF/4loRGxv9nqawgsYAk93TV38V4Ln2Txvyhki7XDQe/nw+gjutdtt1z
lbFD1hTON6/Z9ZqAITjPQkBFUfu/o8dK/waQz1Oc3X20ApEU8qSdDM8NVHhdt3leY13Nx5lkBebC
obCkmD2CMik6kScQoZGCdtXUKWOpjgUruFQMHSmJTLR62vnNFuluTbTiSmkkUwx2l76vAIL5UMPv
k2/UP57ylVkQ34dIMcDlcro/gTUKwqsV3AsSENOY1ES3V+irPVsPIrOBai5jpxQKCsCKxhRoccz3
qGLEI4RI0pQ7fuaFC47TfeU5JzZzPANXe1Og/SOV3W18DyTAgEogDGMiAAQ74nk9bAn3nZILuen5
RUouozuLCm+j8TbsjtjWDTLuJJsipaV9WaJ7vxObwqNPzkR6CBNIIXUwaK0o2ZWjDg8z+pbDf6AY
RDFWc9o4yDFDEVxoPlci0dg29PHdLWzx0jCMvr5kC4tvCzvYnB69BS9XHeHM5WobSTNsNNHvbTtY
4C1a/AWcpaqXY96xYrrJcAVdr7tia04nd018VwSZOn7I1/Ty2CZuZiCBKxJgAVCvbL5v7LjMAgES
gDmm5QeCCOsuM1Ed3cxXtAiBLLSWGIpSHD0pES45CYRBpQZ+P9q7To5q7Jwcp3HkIqhhIi6RuIQH
QXxyR+3i0gtTa4Ia/YhyheWb+qjHbes2N4/bkZTTirpvrwy8G/0OxdMBvn2B3HMiONq9HHxs8Sx1
iJyYhLueXHH+jpCcOfY5mxas9ldprwfuYLaLh1NIJJeQTllq+ixUHaH3PUqzD/9FfGyUKcbj6LEc
K0J8PSOKHtP1mvCcggmYgEKxB1BnNV3+uRkei9fvQ7j8fHm8Npm3MmdfIvewPoYPUMG7HxnVJUX9
skQQKAkmm0j6sAA7Pj/OFlHsIRgnCD58NLK0TGZ2Trod/71Sd7MQqytLw/8gtCW3mq+p9ur/Ow4t
m28EuSZHG4t3Db8iQVCuKYd5lAmVRoCIoKOYJOW5oYOJcgivDUFaCxN4cEyIVFx1/WPR8DadsptH
2r4hblOfNKfW1l1P+YLVj053GEIwOHGnNQQzHLeH6kgkC7/WI2i4i9U7P0N5s/mREcAkK+mpa3Qn
y0HWlYan/V6k1ULMWyRu0Avw4ypYkWOWKNQOWuyB5NVLsZnkEScLmgNNFXpDVjylZNhYzwtFX2u7
VCzcfnd6iPHDhRHr/M71lxP8DZfUvWfNtQ4hAE6ow/B/FF0X9W2mi6JQEV3iEUOxS4arnga3l7JP
Q8QjlAJmyFHcDgULdVT99jKmsi1Av9kOtdab9hYonGCrLywYUnfvL3QZ3wJY6mkrmNeL3zd1VIIG
r4/Bnx8D7xagLgHSEtYtbzNmtD4bkGuaN4Ld6Eof0Xmctpzuy9W5G3aDChYDWgbOPZozPoNBhAwt
PEBMMDipN+5ygbl/AYFfX5NpEh5wt/nKlrBNgdYVG4j5cDs8TMultrvqNYJJTkTF7pWzKwUpoHfK
ryLoFuWmkeJuE5+B+IGDRK/frNPknr09SLwTuxGSD+ivbEe7aelzKSC4JkSTga9LT+rpkBMuPswK
PFy5B9UouT1XJltEIc7KffOa5GcLBlX2OySRtHWDQ+Rf85YGhVU8zJ/uH9KMnnnkzeYyOdKk4a5H
qHOP15XEf0Y4575yBfKiMTTvcaninQUaUYo/WfcPr5mi2MIZJ7t3Qw3zTqbnR3ifoetX0WMZIyhh
s0Mi1mOzimzjxCYGhbbHka8ExILutaMG8Sc1xS0wOS9Cve4f8kVxOKvwftI4F6ZBHxk68ckEovFc
imCta1YMe1hgn2JXVBKByfM0gJDsOnHLBG+C0mT/AKjqbkjBlBPlKKK5C0SXEC923QEBZfjO1x6U
aHQ8/Ud27M7YDwSR1jXV1TRD6E0bChGtP9gfEX8duuBcTIzrZxLt5ZU1ejPy/zvlC0+A8R4qxFwJ
xoVy/z6SoGIht6RRVzFlOT8I9LYsuCzwqckoJczHzrBZakIPpRA5bBxjGWpJCLMWD5k9estxKlob
E33i6z6dHSGqshMPj3azHVV8It8Uwkb5g9MXkLGwn+pAoHgD0HICiklZCdw+8GVZ6m8fhXg8BBlV
iIv3bmjR475nkYH7D+2izuddjOjiBV1jMtYM6Wq77/Yhn+/x6oPKP1u/4GwBkf0AB1GR6TOD2QNT
kKwERI3mZIMbm1Umn2UflYZ+qZejRHt2avFZ8kRc7FDeK1lfZFfPKz4QH7++OrJ7lmGKwLrxunjz
4SW/X5VTzk1KQHCtr7EOdP1jfiOMF+UITuUEjwWnlEzBaiDH/zZokX9oFqT9+xRiW0PhRz/4Wmra
kJaX6BPR0LQZr0qSqly6l0AQNyGZOHqwh+aKULQYyLBkS3WvPKOkrIvfX0f1mbaPmI1em2VqhmbG
G7IPs/8A8K5F047aGAclmDyEXE/0QnQ7ygMlxk5umwb5yxdrlEwRCYQjxkv+AIGoNZT0uw30ZAbR
34GzYC+yrR4fioxDH6GGGV6uxmnYsO1CMdQYpdHr3HuhGqjrMGPlStOvZwHO2WE2H7OHM/5HR6tX
6a/twwAUKGX/aMiX64dZGQASaL1I5+seysnzaC66i9agGKVY435x7BDHEB1+bz6BKLCFuIT6+k6m
iF0qLZ2VJMStib0KVtJnO2KUJZx88lInCGrEV1AOJPAqo/9xmRUcycf8KrD9MB0DHDoC94A3tDfK
oAhNqPqUqyS9Bqjow+9klEM5ChB+i2jShoU7cggu0MNG/65WGRxGuvffi08yDVVpZrQF9JewdWlk
aydFdKZHcgP/CdPcuOSMJIPNv1PhcGHk7cQpKd2xWCmxZbooapbwhgLz8mMIe+kl77NaIhPUxFJD
vMg3pZ/Fqo6Uzi5iRarOez/sbmIf0SYjmFQTj4t4VFkCaYGdj82Mi8xBCSlA5ziiUIXtztg5o5bi
tZMrMSEPuygucUKVPDrZHStk08iBJ4akjx68gsjlL95Z1g1+u0d6jbcVfZoLAROx42UQm4gxlFrz
ZRVHAm6AClcSwUNJLYUi+YvRKnVU3KFN8+cGUgPSohg6jBi888NdlQS2O+1Vat9GbUq5fB+22kgk
A1DhUofOR42hzJV3pForON6r14Nz7aFITWnAKXAPCcozY6OZ3ICOl+0sGSTZRU5q8V6A750KBal3
069nSARAAy1puJrmcKnk60GfidIwDI+hYx8tzMBv+sQd2Rdw5UY799qGaWxCzU/F1eCCbvZlWti6
2/Y4ucAdFXmDLqt3AsztP8TPSUUnz7im4EcE8MOseqFRsI9o+AlJ+l/D1Jt7s4qq3HRWJriBhmjI
rrbDrZ8oM5IXAGzarbi7roPiNxtLAxYQliBDy1QQS2KywUk0e5R3QnwbGysQ+H1l4KTh5a7ZcIT3
FB+9HWwUP/QqKvB8IdOquXfjIKwizdHIdLHf8O39VV/8g5yxHBgVJtTVy3B0MRMB+V72jZxbyPAg
49P9rKUat9deylNrqodJj2suGB8tPo87BSdP6iE+VSeWWn89grslgJqrxpr6hSb7XULYQmIGLvO0
xJA0avLm8nza2NLOtAc2EhSK4XmOyEpHvN3qimZCVWrxRfzZlRxa/rEiZCXBzXRhNp7WNlHS4Ax6
Hj7GdCU1sG6Bm9nsAzqXS0ykfzW6pezkhR5eB6BOXrnz4awBf7g9pzD10dtVy2pykqmDUmGrE127
xSVYNzNJWSiSTzMt3+ZO0vu+/xdvGrOVT3T/g6lteJNasVbGarEcrJ3UkW24oNQE1rnoBBrLOxRJ
HPU/xCst2LREU5DQg5rOnpPNPDzo5croi5jNHtC5C1ied/0IaUZDejOl7Hwx2Sbo6dsvGaDSAuzG
Qb7yx7mfbhqDXFk10IjbN7gyapOuwZEao/FYewzEAxBqSTXPhf3tNrCtf5DRIykU+xsBrJzAS/t6
9fpeWCqTe7xrMwjZO+gcQNtfFXeafOEq/Ed7JfGJwXdEJKxfJQXaTKIJ7/l0BFV5GMAV1tId89En
iwb6lr41Zl9mW0hDG699bQ6h+KoZp/0ABnu/1kf//7jIdi8EQlALoEpyk2zY02Qo1ln4wHiaKTf5
QqgRlYSc0Ne9HeEEcwZViKb51BmI4DEm4t+/MIhRpvTtIuNq+McHUv0V8W+3Qbjy0MkqVORCWMK4
udhO8N1q0CW1SxOrX/00Mtwt89OeLEwIv1NczyLXl/8B8+fMGduO2yUpfNWHFbF/3kkim/Pl3jfb
4fTiITQLPpBrpQFCd5NQ3HpM9Mn4574IGhjS/jak7gFDOzWn+Z48aVSBWV/ptjdhWshgZFdCFLvX
NWRPJHTGrEDkFLzZq4WJV8JWLU7vP4mMt6skHFmEX3pBIA3UD7ToEEqo1a1RU1o6aWr6mVrNLP6D
Tz2hwkkhza2u6J7PVw4pij4eBw2ZGGYaZz7QvrXvHWlsGmOlhWD58Z8DMY0wOMcm5u/Yn6RvlecG
grTxCGcqeADGvim+bOK6I4saY+nd3jFay4btqdZyLCAGNk7LeQlGv1clPRp0zz8A96XaDKtIcvqm
/hRPRd5z8ccPJQ+28PR4z6JracyhUyb0YVJ/7iYB2wuCa5Rf6qS3fH3LNJltOpd63ObiPJP1YnG7
5Eklb4iLWCdX67hpaY+9iMJdRhTKuW7A0dgldeGIVKKePqZzaSpxL3fKQA2Txi6RhwZs9qbXrnfG
oAFFxD6EB/SfdJ57gdBBcKER269WHIs7qLORDATIOYoGe/6OzogXig0Uom2QlO19Od9hANsIslRa
2ukWB5ByWWW3OSXW/rj2hIg7I61tsz8u/MLhmSMTQGoZ8RFIYsU3STziFLVlNcl7I553JS+LMPUo
xaIRJmsYKUSI3XGFSqkY5iIDv5neNrkOFFlGfMcefoc3IMVDJwB1+zC13dh877vQ92F36L/LtACM
uRKG90cfeIjLxmLSF3OlBnGCWi/JJKZ5RI4qA39awu2bkC09laQ3X2jkCA6D/7EYEynSTiKbL+P7
ng7QlmYFNN0urvT4yIBO7ZUNG4vzAHasgA1kMhXyqjA62xJoBqFSfvuE/iKxkCvGpTF81NoognzS
rO+aOH77IAvNthx7xGFFA6osX7A4QD55lC99ZT9uBgAevERxwKv5ohdFGXtZFyiBFFCUt+V7E9u6
blMIa97QEWuD74DQfkDPeo0DrttD2MdZMiwWGUrbvX53yxZ1sUiyOBAmoUPkwEOTL+ccvQFdywe0
sJoUcYNxnqXuncQ/axZIblxM0AfPQhfP/y+Z2zE/KGugDnEgRJbGhVPR+suFYZQZzp5uwAlHn1ne
ACJgJDhBBu84aNwBYy3drg99KBevBNI4Yql3azlEDOgmzLH0GsDYp8T6Qo263tKDziOHxbq4iIi5
GhI1KOPkmnGannF3b0pypItAXMsefNT8Vltt4t9kesC9+5PEwOFqD9PQFH/3uy3W4na2DN4MfROL
/U0M86yYcKnciiOC7ONElhLlAeUfePbM/u3pBXYgPTymFxL2/eWqvl27rZgvWpyDO21uXrdMo885
ru5NGd06Cz+ZVbI37gz5MULLsAGWKu0AFSRmNhvSGgIf4UKw2clYRrAaepK4qqWalv4PxZf34aAh
oylBU0I1oMPUQooOsFCOoOSikZ2Z2VLf0gltlb4L6qJtOVs/QeYM61vAkshdjATNeaRezC4mfEoR
+H9zZ35xTbie2jkwWMjcEJFA/RolR0DsLeXNE/KvJtUccEXVXBgq21yWHDPitx5pW6F+UTTkWhL0
l1LIQTT90QvVFDtpCkZPLesOz2mNZmD3FXWDnOr+AhSOrdDWW/IF0etjE4r366iSP1KtSyozleey
/ZPEmJxPuIYQVWtGhsCCXQrlVa3x2piQtdv6Axuj/Jhb5MUwbzC2pYpzU/4MBLH15HVQXgSdjfYX
068L/RR5GI3D/UcBX9S3r5srm+mmLMzTqGmspEn1nrA0H5rDWUVOQHNY4n4+CJiABdhlHNo966wx
Y5hndzPg88fQ830vVgrRC/5c5bEZrUi0Q7YOhIl21MbQ1e7tAaI/SsKU8bi+OhXAZsXfN9PEGKk2
7ZW/FH73Iv9i0RTGjTnhQqy4SwPlVCvhlFa5IJ2KBInyDOvezOOwqeGo7ovum0gb3UwVq6EZSX3N
wcV3ifESC+TfAgQ65k88f/zXtmOpbFESs+q8qVzEmo+lrdvEnQnbsFiPzDycBvAQVXq+XrWv5GmE
ZWauQwI0djolkE0AzdxgvT+WuRp1y99MDD0uh4E5lFBeZ3LTUKBBG9JCNlYdEfXrkkjbCZogFn7j
mohUmRhgfnOdRv8qnPWvcj+NdgVyQ9Wh+TLZkivJRXue8xfipfi3gdlKJlpsbb07pKVySWXor8vD
Xtw4szYPEly8ex2dcB719N7nyYUcztIYXjVwNI/EgxD3Ht4DyMQigq5QBjDXy7kx+NA0oPapJORk
3ykMQdc9+mwceOoGD6AnznRKWEgsfTwbvanTuOBPtdQVYepFhWgju+KOj/2QFfea83h/KXMqW6EM
AqwmWtTLPQR4K3D0q0VxSulvY87SLLJVEiiIQnDW03xSoWgzh2L4afB6tQfQLhPVcXm2Wnv9HjEP
C7ln5dHuBuGxepxRvrLK19xx17nbB5h3pDErcZ1Rf5BjZQnB62Vtf7YCpl9Ko06v1dnxw6o88aVk
8R0xSfyZF+gR805d1JLVFFzpD4SmB96pa1bE2DfffGScZQ5ELQ4HxRwHwNc22Tx19GVesxw7iJ7M
/VBHKW4ps/wzTU+jxenpjHDZk5tdaC+zd1uj9JabiiHFENM/BMKX6C7YK8F9lMFQvoi133IcXIAp
7th1hBCjyG9u36+tsQqUSy75tdEzlsUe1NUjHvRexrMOzHAVHfZKn7J0chYgVqrsrUhY2gbiYYNc
fmogobAGKUx5d+LoOGWDT9re7nC5LN/vKWfUYOMonvUL4Ak+3Q8lMJWO2sncdOZkU0qKqIJ7MaIC
RW7V0MRNX1w9u+oPwEcmOR2DEhNw1n2W3UqdxMfl33mf/Etyo6p6nYnYTJdZHk8ka6irmxUEyeWL
IsnQcLBpodJUumnvpvdPy1MAlP8lvn6K4jvtAl2IFPC/LOK/FUCtig5FCjkK2OfK63cprhDuJ25K
UyNPxKp46uFG6NnKotYdeZE1SB+MVE7HoWRFU/izcljKSkoDTzoCVdvBHp+9Zoa+trG84bN8627L
YbqaSL4B9WnbdLS9QWhD7BsYMeFvH1YdouVedzuSEQ2Ygx8J875+WtF4aFtPl5SiB45A1SyOIm3C
qAbP2Bnq4C6tV0FF4JOtcx+ksXC67QYGkItU4mhpwtDXoemGPvyFBpVzX1PkYniDvN6XvdQBO6x6
XYAZjlad65lrC7+WA7IP44+Am2bxmZ3J86DNnEfvPaAJX99ZIiK1t+jKy/aTAs+mO36wlNBzg+ri
7mmV/aFPK40rpHNp1urbqLIlMCU4Ud0xdjC28MPVSJny4Zrfw2rVrPlj0VxDiVcakkoFi+TjibVf
lbtR3sYVermKv2iNX5xGWX4asYhxTQ6RB5VEzGTjUEmHNiiV5wX3g+gmENlLopCcLtgG855QRs03
enbzcvkVZAymuHboHIL36qHJU5NMaBOk4/33XOSeNlX9TVArqAv76RELOVbMU8kjlWzx5juHowcQ
aliiFqGv1lto5RweTOgK7IK4B/OnqY4C4bDlnOzzec2y0wGrBGz3tlKliuSVSn+iGf1h+xltmfxE
K+dZdKHNRtVQHv4ivr/GO4suyQHC4JKsvLTnVGxb6FiNZUEnAtQuHRcb5M8ikSwrxoimSLTybLkK
KTCvn7ysTgh+pQK1dyYB7su2fdpDgIUReb6jQVeiyAkTHWzzfuSC2BAvFHiDabAJ1sBMZn7n9/aq
DyCmX6lh6VPt4zVSLamfOr/nOJPeCE81pfhtfJPYyo7yILab6DouY76c1i4oimdE6OOlirtxTLq8
zoxsAWDjj0TFjQM+8GV/PvGL57c2vq3C8kILq9h/Id96ugJ4e4Udn8YHx+C0zt/L5u6qwz+VZef6
AiBUMGUMpSZEQYQMO+I+MF4tJhLrdAxIwV+DO8TVQ2LvrA0MwPAAS/rSSKuFGl+o5rCqYKkAidbA
gHYXAXS6H+zejRJF33dIu4PpRcojIynYdVeZMkvSMSy5b5WC67Z1bCn17G4GK5uKH00S6FyTeDti
7mnjsbdRTLSNR95ONF/kFv9UN1kK7ezYCbgqj2aTEXchBZ6UkWglJU8mTgw3Xb6mmcPUia06q10B
aBgA6th80iQvyBG6N78lyDSTERBpka99RcU4fKfHUrJZJjZIFxFhrOKpRMxo6OGzMfW/rmlR9vQf
3aQ0VOY762VQmgiaGwjTefcqy39eTFUDVmH5BSKMwoVa+GztVSshC5njW282K1jC730E2TVtnl1/
iWXzFHfpPjCwaHPhDWXgZy53VDNeZJuMPnmq2fkkJKcn/n7L6IeCVfeGxSR3zGPG/h5GYMVO6z+Z
/89HTxaNZpdcyFpT5LRFvGA4d1aQJ3PF21At7gdApSS8OaHjY9K/vAqunwtjTJezbpyy2+fS1DB7
JzUHzzmyrJqFd/8CBY3cPMLpxYKgBQ6mRJ7qbbYvUTFgwY27YriLcHK6ItKEL04/R6f9uENEg+O9
4UFTnqcIyIxUjqF29iLoC4O4+szjW75E5OUDzIEruXYP336U2+sc1KW6AcWqM9Kt6W9QuhgHk3gX
CtoLmqmoQ0UVRsBgbP/VzYobf816QpuM8uyvRqoFXhynMkJGpGBYEy2S6J9tzAsjCjTK82hzXvj9
UOrANYVXCe7GB/fdjChNOCaJ7uHfZL0QVSnUZJz3ihjTZwyy8IF5c6RekbXJWAWFLJPrCC76d+tA
4pKlenaDZeGypyPPM9L19L9li3stN2dE7d8S1tBltPVZMjxAx7pLjV6qLmxToyaFJCibDBTPwA9m
WHrhmPB6DUYizZuVpI53wSy3vTdonS+nBC8Riaw4sL4a9XQTLiVXtHeQTnYSqNSVSuiiAEM73zvO
1yeTw+xOAe77LOPyNymsJKhYfKtJUctL/kNWePJP8qiXfkyd5CP3PPYsQQ2GhlfYJhnQlf5Yb1xz
Iyic+plfESiMEU7uQc6Z9jRsfwojZ9TY+i5qeJ/HoplgA+7m+ECnRMeEZyDUefXc6dnORYzhSu3e
az38368fxl5aspGBfrSXQJBmqGaCMen12cZfZ/33/wl7y4OkEElCjZaMW84Hl2zGZ23kj7Ki/C/b
NSZLEb8TKG8ZOy4O7jd1QrOsFl+oRV7cqdvjtw66PX3xmHrD/NdESkowXmu+B5Fyx/sgy2gl/+ao
oeEfIzhUlCRnu624UORy7lzBxI+AZoQYRKLoWay3CUZ64553lwaeGSKtUa0+KQ181+vJSy5CpTxF
/YiowvloNbEnpeynvo6jkTs+O0dAQv5zrFJIVjBR2DMyjjR9tNHDed0vj0SvXVmEpCWM+qGXIY29
fEF3VyhmMUOvjKMVDuMJy/kZooClcKZILbrwgv/CDK1rPlAJhERdGkpp2ru3wQS6g2MyK50leSnH
46+O4OHnGhScs1wXPazv43G4QJTs1RbLXWcPPhhbHJaX9gYPTEvrn89qzckM9NAist7del8KQcdx
bZrhQC0yIPq1y7eQvIlu8hd/ieszIsqJew5UDRjkjMTtT51y3ry9J4qQHwA8Id2kxO5qJuxD+cmo
TAlXhufBgl7jrjhsNwksdZs2QZvdYRRpkepDsrxVtpp+XDgcAV0wsw/LWTjrDTkMyVmTZCdLe3f6
eoLp9eIpmIH/Jx22mx448BUWenJpQ4ohkmqHzPHzV0cyTzXqVc3b/JekW0jyE+Q+qfjZHf1cx2gW
MBLzGZA8VV07YlUTzK7w0Cbxa0W3t/IR+XpjquTKFC60PeaTRiT6be0mzmPZaxKO+VUQjRmMyQGr
Bww9IHEZ7Dcsk8fRovT4zf9zGFLhv8LwNXtQwemP8tq6yBn73D1Ol2MINyVV7GSfQEF2z5WC4WCY
d+vh74BI/syz7aeS6LV25bFiM09BfUUUfisVijxGFGcoyVMcvHxbuHCO8BKRhKLEqY+VLKmAvMnT
9l7+Y3laugjr8iUC9mkkls3kqkJdEJfQVGVwF+hKRYAmYUHvie0H8G49XCrPicMS8pMW2xmgj2TO
kgNoIlprEzQPHGoBReiM5C4nDcmuzH1LsKKWQU+PwCaVE4GgeDZMSkBXbcfF42rjhJg9F+jZXrFT
31M5YIi67VS9rQ3KOlVX0d4h7l1K9S+YT2W/qhCmVwC7DlAhea2wbpPVvhY54GczWiWpmZuPoknb
ICNCNjJDasdeKqCvt3ZE/cturLDqdKCXIOepba8/Fr9H+arH/Fp9eXPG9F0uBX27ni7mBUrxKzRD
8l3GOPICraR0ki1RAwG33OzyRYUcjU8eKK3EzXgjtMSRatN7Ws4S0a9wYdnblhLy8za6+vIJ6iXU
cio2bBaix8DWNQRcGlLgPLnZ2ZuKeYDTOcpahtpUrY2I6yfreueB+f9vq5NOFWotPy0DtCNr38J1
C4G+Nc++9HmS1i8No7SI6DTwAIW1z+Wq0XtTn4Fgw7jFAwIb2oe0Jwu0cXg1fTIXFYgrB09Qy9HQ
3RaEhlR0sWjI66hq+HFhnpvURJp4Z892qZeaurskUuI+HVPjZfutB9wNeoAycrLxU8+2g8NDr3jO
5QLThiEQjzhkSMp1de6fTjgm7OrJcvo54gMQDGrJGLzAs4tYzlzCHHWPo3LIyJhHuEwZox5JbNNB
YRy7yHa/uGYELladkfqp0ELSXIczc3H5gulK4nbC1KHzZSntjnjsBrTvMcwm1eeva5oiCrvCGJbW
ez/gncjADxBKS4WXWh8gTENbbm6t6XUuvnn44eeeozDCkY8RZuu2HQDvxnFch/6PZmcPdQxW78tv
aN8lmly4rhGFsuaEMN8y0aLx/v6sKGHtZ02FAdsCmSbsvBf4syGUPPFwgDgN2On+lsd95xNIr8p7
AF3jGhheUXbrttr10jeX0lIdmJ7Rn9GWiUqBfxpaZludHwz3zdJcICR7Zahw762ZTzwm4jnZtORP
DHcprCTsmJDefh3jA8ZWW2OMoZdsMwS2Kqf961nj5g9G7UzpEF8D3CkvwoAs6yJ+HFhyG9KT5VhI
EZMd7yk1OSHdcQQuCeat7iSbYT97qZOxWSGSbw5L2kxAEYuAMjpz4065mmAr5MPvO8LtrcP7raNU
amSgiZ5SX1+3d3WwXAMHfX07Kgw7hF0H9PB9YD6FrFaVx9p2dtK6umkF3BOhl9EjW9w/SDOGCcmj
fnuxFEGkAFEZLU/0LwkaD4PNm6Yk1qoKGZFbGKPTJW1/crMnpPrnUjoonkeIPp85f7WmjJ/wz7tl
uRsxW89Eqiwh4GNkyJ6/OfmlfTVROpjyv5JrVfb1zB61dckIitJd5/BA44R6cwLZVfbFKl/qmuc+
W4DvXc1nFSUi+AAUkeCZQmzideGvLAhGdrZcyzYsDPD5prxAUgVIuA+8d1Tbh6vz10AvLOGAXUL8
N+lDcNET78jC+MhuWg2DEmae740vmTkZhqEQBXa8c/yZ/qKZzDIQrHEJ/dy+Dl2LFjUQtJfo4p0T
x2n2iV4qrajhRpZdbCRe/X2/kV7D5l2BqsZ2P+DtbHAcxTaSpv2dG2j8xTpdzYE+hA0DXpk42OL7
O7VQGuWr0eOGJw1LQwAubyLn4o/izTKQJVq1nqa2WT1aExcx797MWK6546mYNsySHgMQpyPAgBvT
7WUcIbsTIB5E5BO7meziXrc1R8pBW7qQq0LIm+TcenlI2sTnSpb0d/3h+oKLZ+QIgoPeZ4uARlPN
gNgI+Wf091GL1BknYZxg+oPlhN3GUlpjmnT7EXopli342GUTzhkhpK0VmlTWkgGB29RL2HCzsv6y
NJ+YGr8irTsA5wnWNQkqoQMlsouD3iDhefhMOP9uAdN+rXTgWhqtCD+NIOkhOVbLNPiDxBqHh60R
F7dJZmAn1zwGjsvj3o1Sq3hvGf1bZgd6snpxL0+kBZ6uz9h5R/0YR5vuUd1ithI705YmGPRYFXDV
QmJkVBjFTCcybGFnY6ATtzTeecppskWAy7EgNmhAmomA9MviNdghSIhmk97uhArNc2wY38fYHf5D
4m0qDWfdauadPrxEfT0o6RJs5y5Pp2xtuW8binyxazMRCm4a3fw1J96thcmZT4V8QUdrb4A1bjjM
qemleiXQQuDYUCioW+HNwoJWj5UjlIJM+JSfxFjK7qgz1nR0dL+tq0ufC/Yywy7hSw9sKoVvaRI3
0y2OV8E88uRs1X4tMdIje6csBBN19eT3oWOWiVDtjgui1tYL4ssS0mxAxhkDSFSeePTofxAaHhBz
OFjYUZwlvXJ9v4AWpneWugcVarD++6Jbx3MGH7JKq+nAzdQF6wXZvYjXMKMjHf5nDIP7J4BzZEiE
Rsd6M5RFlOFy1WoeLlWlmo5kd0pj5FFDIi3+f1DRFi7N2baOmTejB9T/hb6gViC1qcqZPMDoI1jP
XdkuxexX6o98oKWfrizhrHuEusXfsPhw7QqnPExJMyHgDitI9rmpqPCMgmAc8kpZR04NT5tjhMNL
ZqvIh/3Wx6yVb6k9HAepIoOf1YdrMRtZcXgcz62i14VRp7YTOWcWWd58hMJMiT/VZWuD58CtUcKJ
Sd3P6a8B3uFRDze7Wymy8QDfcBR/Dhifn61Rlic2Srgd7/ssk6X2/sGnBtn6N3tstRkavpRBtlwC
c+i/wsTwZG8xCnVCSQwD+Aqei9EBbwKhKFvvhmNqZRptomPiac0PHgqE9wAiZEz+KK1nTa6I6BNr
DuAdE1OKBOipIR/wpO4qXNEmoosMppiiebUdBYAmONZqB5NqYLalLY96MQpT/+HkrD3jJhAB+pgS
CzJcdECh6KJFaBapOY0EoAMiyDOUocae+iic/6e9fXqJ/a6FsIBgYTzJUw0uRMiRNDOBPi0857zo
hhMlcK6g3TTSrq9VRTE8bciAHR0qx+KHhWuopv7P8jvh6vIqhnrTGJVGaL772bQstzxe0sSpdjuo
aHMwFOF7uKWwYTnFNN/3B9oQfvQaU7voBBMbAWM+7utxSPuh0DYiCcWwRU5L8CmpYvuokvbBdtbu
Fz+9q0OorGY4Z7w/jXgprwzxeZly6BrfJXHxWH7iloegX20vNU3BlOFrdSLCHWvt7DTuBeaukJgZ
2XUoJsuKGYSfIm8eiEq6JRFNPGJT7JG2mnjG+dUJAZBHzsWCW+JVBtgyA1JFW08u2BAACTPzrrKI
ZIS24VUmpTohXf5NMASyxU89FiwIRnb2lK6q0NMsbbm0zptn15Hn7tilkG6DcAzwgc6Y2F7Do3st
xS1Lqrdu3nlNArLlTCw9RPpvRcThGUW5IX2dhLr7TAERtPj0IZDvF37cqpT7114iXI/1rNI+gA6/
kqYupyjAXz/09MTIbZ9En5LwCOzvGc/tEeqgXPGEoQkITdWv84iRF4QdX63ACNkqp+JpXIn9wqKF
K5FddOz1MxAmZYCErrLCpsvibEL4+EFF7K2lsYs793edjGJdoBfTN0F1SFMUjAF8FF4wbxZBnnKI
A+SdfWFJ5gAI3F/OkMJBXcBYDyvjqpoPxJYYGtY5W7Pgl4NgKxAsPgdtbw+y8JXHuH5VhtgMmf7r
HjF1TVxJLzdo3QxpyeqrDOqyeOlc669wZmlIUo7HHmCmo14btPWh4BalvHZWjXGg++M5vT6Fa8Iu
/z+6Bf4srMxLVPctOBjiuucZt0l21zpqgboyvVMOiJsT6EfEfHOL+cgdCi02p62CYPq5Dw9C+NtD
rYDT3Ke1xMN8ftO/JsLNrn4chsoHRHhRXRRzv5S2Y8WZ97bAPCzqaw/n3zz3CAaCiAHj/zSizwdv
rE9BGHIfQOe9Mgp9fi40lGG1F0OccSOJ3lTTPzekwa6XzDMTIOhEKjYV3/rmmlU3fhGWcv8DbW6p
anPQGBZIeEqj5dUNTZhq8MjU2FLKLqpKWNOpsId1fhCx5XcXL3RnJ9sgVg6EeOig8WW5u2Ep39hg
KdYL7DDbDz5hEQDLdmbH80f5p8ZD+jBdAvwUNulcF1vseRsC9EOSThdnu1/rzmWZ5tOakKw8pBFE
Nwc4wlnIalTL2XKDF+Px6+/mCnxXr/nlRTYTRafusgprAqPOOpGWxqna+C+l2HPedKngBATnCTte
TniMwkEpsgFEepHIfOXHiToDUC/85j1ASL1NCpHnhrVcQn5F8M+/RJXse/UVcqATD/pxrbO+aHJz
4YxzXlFPUvRzqT0Bed0pXbGWPfPTybDcS8cAdgp54iPnKapBbsQ0o9gBJ9ul5QQ0AgtvhLJq/HY5
KK7TRDsgu7Wy2T5MFYAYfpKoeoei2cC/vKTmT+18OhMlfYMcBeEauO+Oqdcfz225RNKN1dguyGm3
uZmi9LZqOkGVlWquFTl6XYmeku4srJzYD5GcAiQTws2/eHAeUfEn+JcIv+iMusUH8DF93zrNORDi
+ZrRS4PaQ7+AAFO83jQiqV+8+i6EcfMmkQXJ9JnQeOqK7WHlKvrYnZNm8jV1bjYTfsRfdHxoNzUy
dDbF59zIdLS6GECtDJdzLWqvt0rx79PiaP0snS/lnubzx6hSQl0c0th8YioTQPeX91l0aSKJUF2s
3TyF/apactxx+HydXZTBMdkByrdmJruSiUW/3is1uLEvKELlmdYmmbqKCTIpJIG3a9+rj+P75YKg
4+eSgUWQ0pm/I2onXXwzIwFCDdBFuTgbar8U0HvJozUMGWeoRVnhv77mQ5gM5fXlQshYcPj9agbR
iCWXH2jFkS/A0qAwu8+HeGe4hpJPCk6ESk2zDvfurR4Ztgwj3snCeKMYDi84b1rtqSNv5bbMV96Q
z0B9GhLP4E+WjzW/6e8j0QWOsJAMQDpx/2anhccWKzZjWEDnezZM4zA79UdjlT4cz9qDAxuY1Ua2
2hHL+kY+armbgtOxXYMWX/5JBYtVUrHV0QNKoiW2nzcOsFNSiXCiC48kVfDKj3iOQZSE4/MXODcq
kxDBhHc6+hpp6r708a9fsGHNsZxsh5yC65POWD9r8KuuFD+vbx063OSON2hpsh5Xv41Kn8iPsf4p
JrbtNDAS3bMfxofHyHipl0eZV4hQZAPLdOqPI/GjjR1OcjayvoRL4JEGbFbNO2LjNKVaZDe9EfN7
6wxQxTZdAXLvXiYcYx7q9+sx1HOeQQsCUrrpgWg91ILzlGHmsU8ihB3EkvttYNwDerDp1gqEjRDW
2UEdHoLG/fjl5jBMycx6toLaX8DvYNy4LzmOlMxg9TO3meUqQn+ohvNiQa/TyntODUgCbIu8X+1y
DuaRfBqM4VrnxHWzXBCJzdJEzXHpva5DOKjv7DRoisuOAGU4fsqdVV/kGsqZBveuFTEszOl5jDRa
Cgh8Y3EThdI6q4P8h9g+d8Knfb+iCjTn+dl6KGJ18o8oseh3PEF5pLg9FIM+L633+tmNf2K9/foh
Gc16+u8hMj9nYuqDJBgfoOrm49hWf0qEB7f7HEJSn/hpHCJZDBUR8MiPV+xyP9X8yShTyGfRbMtK
udoMNZZtTf7EtqrIFTbny6CyKxQ4BnviNe6E0FGymIhsDuXMYDrl7asyCL6wokc/UzJPM9na4aNc
vnyg1/JsexAwLero0fp2mdlZm8HyhZzHmqCCMOUBuTqgVLIEGvG+lFaVsGbx5b3uHihcdC26vUuh
wsnPtwEJfgv+UvMa5IY7stKUeYaCj/ebHs8wYOg8yT2RxK6kdZkOgsMJkavIVXRZ6V18/3g0H8YA
x6MP2ofY47OPRVEfuCQNRwN8Sm3pWlseKBhlKxv58PvU8fOhoVH/5ugMtTFwudQWEwGDAiFn7Gug
XZxfn32Vt7LJhNTDUjzSj4AARktVMmJJZX+5fvqo1I8koncix66n6dJdoULfKCrkz7kJ2nW31oe1
zY2R72LWAostW/ydE4PYE0+Ce0xUmm/Y2sB2dhZ9UoOOAm3qI1iM74ZS5kegpXhoNK2zK6LwYfXA
Wk7yBl8orin3l5DTn2vDf6vg1D2PqRX1PRO/FEhxNQX1SQ1FNa3iomEs7W6JqriW7Rxqd7S4JvaP
QEmntfr5/RV2Me3+jiJ+U4NSVlK9HrAzGcmlLxYfgNb7SHMdzwueUxBdctOwlzbrzLMsaHUcrIyU
xzR/MZvjVE5wfYHaYBv57+VJAj7kQ/kIsPDDQdLoshY1eRTmEC2YAq2fjzxD6ReR1s9Empg4NA5C
N6Hvz1yr9go8VEsVMBUajnynlQklzFjPtvP1Iq02GJ6M0bc3APbmPR2ki1S8V5ZWWvv2KV9T7PQg
LRPcVQJepBy5rZ23TS85UU/4wsrIXCuPQ5nGFu6F+WH9eeHTp0Ao0kgQzbTkMBCJ7XVYvyOwq4Jh
4gyZXazGb5sklgTA/jrMsles9BBV+LWDJrsslfdOvsA1ao6mektyXn+593RD2uyl+RBc9rwo3p+o
nZkUww7fSpeSK+AgtycI3ptDFMJ4q3iqHBnhiPOPd0SlxT8u7ZhW8QMKcF+plMDDD5Jwb8eHdaRR
VNX7a8YtHCvMBpv2q1S8cJXQoIPMT2A1eS+9wjBpugh50BjhDVqDfmjTP/mr48/YovJ4NHLCvqeO
x+p/qG/1MQjKNu0KMaFv7lqV130XoGlTsxE1ANGLlCQV92IUEzJU0ydE9y+TSfJ7AlpB4frX/hyI
y753VDcj8n0Xjpru35QXPBuMB23W0mar2W1StlYW4ALF2L6PI7crcIQOvgERPxEzlJrw37HjXjVw
27iPJjXR4hLsKQJbkDd0sotPsGpbr/RzA8iaNG+tF8S9IcC7ant6e/rQyPXI+r1TW5CWVQEK3aag
jYqrZ+yJHVU2B3kRI1OjA/IwUL3/zvyig3mXUaB2/a9Vv2tl6dB1KmDtOveimPVrvCtR2Sdya9yS
Xt34AMAYHwQEhgEKp0bZXaUvpJqIg/km1Xy41qEKtANnqbiQblnBUG5GZbfzDLFY6YwU77eetqw5
EjjB4Be4N+Kvaa8cKMiPIfAwG+4Xg3STp2h9ghMmEEVAlpT5ozJd7C047rSh4AN5tAWV5Iun55v7
9pddSirtqeJiqZWJU5suN8FPZuUiITv+N9lAc6md2PvXh1Wtd95LuXvdx4OkIXhmwn0cpfXJAPsW
kQYfFmQstG3VD2rtPOWVXbHukxN3+TZtNUTdqGGn4mc2M3Fj5C45lNSqFP/mU0INYGlfIo/VPUc9
erVk0JqaLqm9V9kOpCF9Seb0XGwPmgGfjXmj1//KjGoTbp7k+9JymAHBuM/y0P/6/E/mgPb9f2Ft
kWFnK2rd5n7SAgX+qjNk/ZdJt8HQAys4CvYe9+9EDS5rcpo//ey8nK5Bg01iHJujpwWq1mV2ZBGg
0QyqwhYO/ap6DZU+4Yeh2cr5hJOcJ4XFpoUo7AoMAaCGpWd0O8T+msioRY318o1J4vocblxD34Ca
rpfcOiPK31HJ4AjRPVY1AiZxm4hn2Baw23UyOYSy/toejszRzrmM7buSj34mwkFvlcNkeT9YBCU1
LFzpImXB81Wyj7YAUgQLVnjubz6lCHL4wHqN2C4TjeT18bQCGI58o679SMXISVRJ7wbbRr8Ku5xL
L45ql3+7dA1ug2/cIFLXWe+XlgPShs1YZaiqxQ/nr5zSmaZFDxtaAliHY+gRPckaolhGvoEIvG22
D5WzEXDxavi07rxBch20Uz8STaW8/so2165fUQaNgFHvOHKwL0Y854zNyhVwjUW8pf2SXwy8XtFw
vsgjHpU6MtQCilij5OchL3NHjBc+aGcYePjUjGn2mXqYkB79rWG0pVclyAVppGiRh5/NXhVp3mFM
v9APQZo+33UEfAs2BfJ4JAmIkW8eg4K8hc8OBdajk4PjH+IwOGaljI5RvjHWWwCs/6dCzYxwG3Tt
loK87LAjhWOK01t7PDsPqEMO7GDRg2+QwAJauMNP8bMucuCHT4Eude+yCXUGkAnKxOAuTzguriir
Qxhja78coysI4seRnOk02qKDgkri3Lz0qzf+ai1MLrH/JSKDlwrNxs1jNjqQvrptEm8I/pWgqO9Y
eGN8Ht7kA13901ptoGBYh/B/3xX5XS5peDEnmQF0RoPZ2d4o5xBA8/ATkjxB7vjL5voaoHJvS/ZB
FYkC12VeXxctM+WkiqDi/0LZFz66TLkHPAQAh7fVajRoGs0iN//RbDYj3V5xPQg854Ks2uU18wuX
ZCqc5cv/mGe/JKI6w7HyMK5r2I1IDavuNLzYZtC2hPDflMPfBeCZej8Ynk1eLmIE2MOZyhgnTxmJ
DsuqII1/3BtDLxlMabG7fB+v/4OEhJKbdgphRG9GaINssaGREfZVpU3yJluISeYGy1B5DzHSLiKR
NRkuZUYRuLEXz7LTNAP6T0JD7QVrVFFAU+TxOkuh21ojQ9huq8gvl3Aa7ZOzLRdqo47qk7/ujoeB
mmfNUo38RTZGGZc78WxVINVsw7RLHX64iJK8FhF2bSEwB5k0xy6NNrRz9KvnvALlAXhIZuXuRbdJ
1fjO52mYkcpXDtXyLQflJ7cuD9X7DBcET9fPLpdev6lnca61azo9wgm7f/+gIaIhh9pGMgi9bgFZ
22FKhorhycZyG+xDuqeoWw0qE6z7NXdRWm6lkbDaKO6ZKhUQzTWdEblc5MxL9sVnc1xtmG3M+M9O
EMkTq8v/oTzqeqIw+YSIJo9a1CxveNTRZwtIojH29BDy5aANlucb7Anf+ZlEj/m6yCVEMz929pi5
phrWZpxdIoem/E2qO0AzwoM63CEZmLnUhvr3bEyl/iQnrxfUSZOrXkUgGWXkvZM/B0zzAR3TTxDz
yv7khS8Ep2/8Debc/Gq+YpGRvD+IeSgXpRAb/YNJdDkwW6yklJ0Np3TCBqhnqUVwVeTkTsQkY6db
hRhnPCGSHE7dkEWDrcxPrdq2p8fEkOTUJiyH2e222BLchvVUuVB4A/yayaYWheoXpB9y127OW1Er
RvFx7566NQqIJBi2n4riT9PQ6ivk6kg2QuABiQ784fNdnOPrQB5uP1TXhh9vQe0VRoj7Hbdja1I6
9a/qkWGs958MyNrnCf2WsXireq6CjfxO/pfmNthjlZxTxHF4//+19HdAp0FdrZD0IW4IzCJUQil0
l3vTkkhlazjxIH7bH8bAMpL71W0MomQNfHNcN0+3SRqhr+SuW7ZCQwXXmu3AdwwpbMOiCRNQakEF
5ew3iDwO4dB07kYJt5eAeHhMh7M9b3YEg2ToTdRCsAdJvpTCv3ML+W4Fur2b9gqs+tYGWqZQagVp
Y3rktjy9vJjMZ94iPu8BrC/xD2MUnmAaOhhQU9KxqdbHQDgQrN6Dn8riMIxNN5uQSNeASQeBOehc
HsVUcSUb1t0aT9yZ97ABOs8NiWpnyULf/SI7wUPDdLbLOSYfeRr+T0Fjjaggmtq0CPfZS8Xz/pDY
tcZCczSEAGUuj+JzSDh/8CSiw/deX9b615Rid7AZV0IxZ5lBxNMcjBXc1iwahubzFHOp3lsJ052w
IK5gVPi/a7rgYKb7UUobalwHdtb0gKVTrRyqOwbA7w2yXO7EewJ29/sdCyZ4dA1KNm6YAt6afwoX
ZvevE9/DqpCBbWPPVM7tLodelDdqKeXNqvNBz7qoHvz22hZrjd5slTUiaJfT8v5kYhfE4UrcQjTz
f/CkqBB4FkoIvdu2G8b5zwnrtAOmoaMScmRKAcc0LxxD8bFNMwqnXtOmjIenSIc+F9Y59pK0vdhG
SS+Y8U2Rx5e5x2PE3QoUvA9wagPhYnduXd1dsgKjcPTVCo/Y1y+kDfuXPHMYG35/fDtebbr3UCq1
OFT/Y5ESOycGdA6ymMiIAs/dxIWIXdNsyKUIGcwdvvNlOJ5Gi6jpdpRJPtsb9ctPUnErV+J1DAm7
3MsJnpkd11kWDS3fx4egyJpdclYm1S7a/IpM7Yru/eUe/RtDdBsv1ee/2ttLg4jrob+ew6EutRNe
Ei/g6cln4SQaYOZxBwCBujawRyifG5YxYGP4rLk5YNU9MQCX0fuj4z1YY1wqYLcpfl3yDNlrSX9O
kmQf09PDiGQC32RyZ7Z7JIMUd7XmHNoIznW1+be3g8oFGvKSt2opUdnYFkyQwUNV27tfHn1vORLd
N37bJQlHGAbx+IhbiXwnZ4BhzVRpHAIMHfhc93sGv+qz19UCT5CKZ34CTq3VjHid8bUXUxAeq+tw
bW/FG2ufbuet6u27Q40r+ydar/ChKSqP7Shonot7ZrO18QjadBOTU/417odIjydjLACoKyJqz2sV
2tXHsCuTez9XvvJLxq1C1zaS1W5Oi2n4Pg8+CL4kZOJTd0VtIy49QUZTWCm+T3MgXKDDsY1xAQfK
0QxYHvbxCT1gv51LAeZeo2cti+UCbGMWXk4fq18bWC569WnuMlEo4BqmylVacrFUB+U35rpWw/rT
N9EMNGF5e3zj71gW0d9j1sx1sfPZkaNq94uvS4iTHjl2URveIYOIlYI7/d722/qRxToMlxRBUaMD
w63im9EGu54V5xnRq/KoyUqjjq2QilbBPsaKVOdhOOz0p30ilLoLhhVGuohoEgW2J7nTqYc1an2L
3Bt23NssMWLk3N4dAxQNuzaUbOvr4/Vi/1MTntHL7m/Oq8OKwWN1I9pVUpae+5moAwrg6jHkAR35
1WUFghxZqYqOIEwg8x3priZ09fhejwK+wucM/fickdqKT78veBtb4a324V5LBGugmJM7RKJureOG
kMDL9js0Ga6KWQMYcH1BHuUFbukHUg9SCrEErhGL2aHh6848p8akRrYGLlj2lPI039WUTr/dc3jq
SFjtsHq3MTKpdzAmKP0u2+ZNiN+EHE9dd5P+OFNKNGR/mpZuE5i/PEm8CQUkd9bzVzra6EfwYoQ3
uH41vp7kY9G7vK1o6BLsq2/r8RgV6iWWDSta+pBm3KQng0H4Pu+3vgIHFO6Uxu6YnxAabkuDd0HW
H7XSFCh5Q8da6eZsfMttkuF+MKLlReYuidk60WdA7SbJdfAwEMRyAfr2Lwuj542j8i+pmAtMcOnq
FkNPPxSbmcR8go+26UdYICqOII98FkTXz7BxW7IiR7atduweoKjKaHCv2DQy4riniWAmQC5mYuj9
bOQGcDj5KFg1XRQYh1XRtkZ5y81qPgxujwoK4/i/tiTu9pNQ2k0v5U+/zid4psczQETuugaomBkl
y8Z0xKO9TFJGD8OB8OKlhmwRIIvfuAvsGwJX7uSnx7LWcgnBasVyfOR2/kxPbEblf0PpHYLLhmkK
6iGA3rTj8i8Egpp+ZBBwCgSmQf/ItjBii/xHD8FcWRhc4eKXFW2TmF9wXJ4koxEV1Yc18GGMH7MF
tpxpNmy4nDhdsi3uGFvZblKzPSUrM3tNr/OdvKgbBMFGYqRLnC3fO5NGuHSqzo+tvCt/U1qsyI78
QJJfxTk93+/1r8fi87Y8wykBCOta3ZZiThsGnU1nwvDKwpn6ZdSWYWU8pLsnlgMYpa05JCPICVCi
YKrOq0w/0xYoj5LcOnK3N1GeVbCbgvG5Fs0Zf1t6/4NU0Q6DOGOKCothE2aQaXsh6nnLEpB75A/l
rqaK/J9bzFAkj7v1HwuZMN0vmkvL0NzO/J7rn/vQyoTt6hLQ/HeuVwy/SzZcXG7UwRjgaZc9uQfq
f1syhfk9w5hRFqrh3Kq9qXHaxuzv+z/MIJ4bll/tR9Fr/YJQV96Rwt77CfaOmBq1JenKrAFRFK65
BkqwRT0sRoKumFoxbnJazHO1V6dKuyEoInCVveiIHWu4+4YyPFRwbbdQRT8XOtlyOnwKrCXPKEPg
orDTISkinbCcQzz/ganSmWwHGgD3/YTTg4WVBGvCr/I8cPMv1yeow+A9SWW96v5prmSZn0R5riLD
tZ5VCYvgB7BCxyy7MpHFLNVHgeCWUHwFEQj21DecWnfgcF1mVF/XMal5jwOFfAbxSuHrevQvSui3
dBa8QjKEabh8qsi+vyTBGNU5azw1ImAUhA0v1k886P35x/oxdAlP0DaSgXS1gehaRXB+F0pv7n5d
PQdeFmed5mAZhDIUqt2FcnzK0hHeHl0tn5G9xMbSl3cDV7ru4JbAmGqXBuYNq/D4HShbHqjcFgvK
C/O4CaCTpktWumt3zDNiutFK+1Y7bgKdGWDCP9iWxtchaJiyeFja68wSdp+mlU1f1I5nQWm3RgNM
QDsZvG06jEafD0Bee7uO8diL7FuUrGYN7pqWfQ27t6o0YwJDwv8XvBqA785Sg4RgUQH46xCxJl0u
E8myUm6C5SMlEKh30+aL80t4hyZPDKz7yaFW/uiuBT0Q+TS0XtWgx5Ig2mTlyvzSsMNW1NaCSi5p
lvRBmLMh2R+2ZdYJlw/z4tz2vS10Ccnewg5OEj3O3EZPaHPumfmn/dPKzGynqfJFEt4F9COqUn8U
VTa9mdgPIJquDhnTu6Yfl1cyaaOlgSaiJG7gX/Pc7CpoWSDR3fOiG1HXVKce/c1L9MqQKN1jDbg2
TlY1ve3eR8mORwkZ7b++kXr/kgu5BotoF8ioWNeC3Gggic5idzkT/rYFBn2E+l1tzzUJwZixTP5J
ceTo+NPi5CoR+dmsOw6mnJmaBCzR2ZS81WNbw3ZLy1xCD4jmM+iPKtJJTy+Hl4VcLmj1kGDnTiBL
7J0gbYwclvRqICl/8Fu4x5Uv0cpXh3Y1+IRwit8annvSNdyTjDAlg9rloHH5N0aohyTverPM7X9M
GaEhxi4GeDFt8RlGrAWL4sFYFHU7kinFGgfXvS7MRYXSy6GRdHpaICcVTENOZuM5j8SG1PkAh0KG
/bJjx3HUxvTN36/SrXt68Ro454HRa2p2AsM341kHfmTNlHlA9ZxrkwlOrkgMqrmseTSDodFJIeTy
+5rq0mPx5MpimMPdqr5AGzak9HL+yttUGdr7DuRMbxJRZY+YxKEPPUkNsbkgexBY7/l1pbMr0EGd
XB3vdxqcincHSiD2g6+TdT3lz7FiMXfaQtvMaszMaaKrTSmMmh94z4LpRQAIQueT2811ulExUAAY
lOJKyfOpR6cG7JaRk/dac/g3uYnw3qmXfdCwJSWRIQ0PXjH5s4xQugsCrxAuk5faZ0+XtLSSmlR7
1oS2skx9UEPlSYxv6tAkrRYcKiM7rBsSXOB8Wnm6kxD2JDD2fUzB9TBSv1kht7ripaDMBwt8cFBZ
x1sA2sjhZ3UorXugWCF2q7A+c4EZq7R94vY8BRR3Fy8EZjtNsMjqCpKCG2y2ULAjz+OEfmwdWYYe
9B+2axY2MiPyqC7sei6O65kC9DObfBL/abgQ/Ks/fX7z2fLwB1dWF3EFA6wsg6M3izfT0e9VjNUt
dFhgEjQbO/KMbZvbsrvRbVlPgr4uEYh4O5EfC9VRQzsOi+08j6PQpHT6z1QTkVTUK7p7D3vt59WY
1bQ32oBdhXfhZVsYPkwU6XgnXeNDMQEWkaSFaVvSCaZv0fBkAGj+rTZsuSBnXDqjdOhO/fUblEtg
iHBe3IFkSCqvO8vQmEI0YZiz0kn91cpfeaYWpaz/t3+I5x3/gyG7kuJC7m/jDgaro+cE4wBl+3Y6
HLN472dLU7CF8BYJMva1k8YHZV+KL1TO3sgvkl+Z7X+YoMzwBHmHrP/XvmcxZMsmVn+50wlAALfP
7/yKHas74SukS5f50j4RUxqww/BUuZasnj4Oauf+2vISiFe5EbZgWA6Z7Y2fdQ1H1FvA4sJ7/FCD
VHfQFmWkYsjJ1m6OQ/K7SRY3vOwJyPWUIaTpOaT4OaKvD+U5izX8dg5leelLJWz6W4DEcxCQPxdI
G2NwxIf/sxuDWPqNoiULlemLPHm7WFFpU88G/PFO5u+ggGIZHUvrykAnB5D4FgYr5nkcNm4UQ/6i
NptFSnltHWJ5+Sj9Wbn6ojQLa95I8LLFgVLIeVEhmgINkPBE1BG7rnoJcs/Q9U+0hrOrWJsA0iLh
Nw/e+zAQoTpTUOJJVDXvL9gsRP8+RZsA3iT1zpYCe7bK9LAHEHH1gSuHJ7U/Nl6s/krOCzy9TGE5
qJpI+w5YXAdKih44+4ZAKofrc8ZPkPPBUGpJrdn3Ex5ak5aT9fycvaS8GgF6w479PGs3wY5G45YG
v/Z1mZQP03fAhH1CGBdi5BTim90uLOxKKHzYr2HvIbGXobYF+EEyBGscCEFUg9I3vj+D0CZFM4jZ
UdT8DPkJnHM0gAASaRDylYezkmGgMmMKn+XXj2EHZSKp6FQseW0t2rrKRVsuYXXQgwXsJoeU22Zs
ciVRVUEW/6m5ETQtt3qi3bRYZElnwTEOl92croEd3FmkK8EJynxx5298BqOBsatE5mqyQ/Kwm9QF
Sr1BLC1f3dwwsWh3GXqR6PhB6asDB76SF7GkH3Ru4svB2FNdvCebVZ43CxWCXFFCDp5pY3GWlkkn
SetEXFPelvjc/8w9GD79jTrru8dRtlNp+lUulVAWmyMseUWsfhrnPW9rmOyUz92ePE4s6fRUra5I
OYbKqvVk03b/WcHcKcjakapIeHHA6kEGqP0VND4bO/85kIIxpnV01+pJx4zTzi/07IO5EOLroePn
EX2NkBo1qlZPsgyonLlY7x8xphmKBMVND6TE1GBNzAB+DxRO9p6hrN6axKkVeHMFpygBo9GF+DXq
mLMvwfiPuuVM+FK/E7qV7DXpM45LSnB9ui4g0c6Cks9sjE5l0XVvIu4iJ17rc2kE5bmLSD5etn6a
Ja2HUVPJu01lB5HAia8qKES+kVhqP9A8Hi6KD5UuJZ6Fy884derZO8iwkY+/E1PhvK2EoEHvkenY
A8rjBlNyyHH4K5fnQoE5GWLfNZjZRnGzcX86tObC7EeGcSHmP0UKXkeE+z0qnzm3pL33KaBYlik2
5gR0WZZ/PrcLr7gJmim4Om+7HKgNJTiBO3UmDtfuVAI07qYe/U6q8NFE74koCrJ7cPtHyzvbjeFy
QaVeM3CmB9nBLFw8k72Yb7eT/tbxvuzdnvqVwANi5IujAHzsTLLp5q6FXVtXGoMi1I7LBy1OX4ch
dNK19w1HH4pil5CQk2zZK0Jm0LmbKT3lNzqq5bFYO987VNw6Ymu3BQaHr9R1O76ZR9kG1W3cbs0G
Xj46CpjqYOwGUdbsKqAYNgP4Z8nFM9/HVEMqbHn4Em+oJTWBizAAnow0nW+v+uTYc48KiSvFVY4I
FTqxUt3WoKG/DOmIfiCRYyHDGtkmdlqyJ8GIIB4/FaXcrgrg4wNLBZ+0GFQgl/4zFxUJLXBJ/2d5
IFDtX5pTNw57Azme+lbtO1Rfkfpx4Y1/yhFHKvslu4GAWftKe9kk4PEDrwC35Ohi3fLEgSSDu5fl
KhFS++a1ATq/qFQr8B3F9aZOuRcK4hAPkc4WOwQXHZvnJJA6E8FQgxceGlLeMgBGSc9XjqD3tDVJ
ohQES9J2es4HK4hdhYrn0SbVtbL2dIsOCFtutb2zseq34o3AxMdpi6pzjYnhfb8rEkERxadjsUXA
OiCAVPvDt/Qsk5OhHK5mq1Xeru/5qKbhJoA4MGf3UUqG3YK7fufR3U1rpA7D7tZ9k2+fS1hrSm54
4XsW75fRUS9ADBR/gKTrvwGtQhoNTJJz7TclQbGb5no++TcvDQu17Gtzqh/aE2SgzNWG4444lSHU
oWbtkygWCe+TMmoF4zfumMrittz6pbTgmJiay2p8f5j5aErOxE3SspQ9UtUay7mxNYft5MPV+LHN
HylN8k/7Gi2w7bv8TKV9IiN2t8gAAak/QcI2DQBhAR0nYU0XxySDrZ0rFEJWKwq0rwaA+WfrH/6C
2D4YhA3ZFcoklABFY87Dtm2McBtz5pbNsZ8DjzGiu19ijTbSqjrryrhygYLbU5GLDD/rfROKUTlZ
8HzUl1W8EiKWkORg71YgXk3j/KDNbMJcLzY/J0FU8Ef4uzoTmyqU8CkPeHqLts8jOxOyNAHeDUCu
QLE5pSr8pb1IDaTmuh0zG1xMl5yldFA6qxnW5FQKcjmPSJDnhqDuS6MDOgQBKH6NnZkcQvojU+nh
FA9JxpgYnoOG01nK2T4PuJJ4HSPe6PzyLA+f1JH59EZVicCFh0yq3cOl48gdswhm1ndYn3gi2HOR
RYTs53tPBowi+ivHbaqD+3AabmE9vzNJcGTfBWoIgWCDk61gDpljk4jRhuN3wbo++HbtaBW1r7ah
0DDvgO7xFSUYTbE3dKP8UcTt5pO4VSoo4bN1TQ2YV9hPZ8zT16IHiJTKv6HYrDZTKKRIsclG5G41
wsP/5etYDf1dBYrwt/nYrezlp16Z4I+ITc6eIj3LbcXFYZQNdTf7tTKrIMeYDqZXed5ov/r81cJ5
S9wKF4bSNh4000dZAzGpiXDgHMhFgmBLoZkG/EPs0KSKQAUisZZpl1AQC0gh2hjw/51TsRjR9dJD
9k5ap/mDyBN/yQMaRtFvnOEfWKsyORX6I+vqDW4+4IKp523HCvZsXANMbe/O2HyvbsMwmemjygBM
rLI+1dgNL7uV+APTuQ9E5llk1BAVIrI1ZhBPpYZ/0R4wJSRd0nxGlhiT42UYKJQRDrvQfkwaaRrf
y+FtvEKbojE3/mm/pq49xoSzmlmTyieSfzXGSUopD9UPVt7/zSW89dekOOMg+mIPg0a92n9Xdh3Y
/1EWRcZ61G5tj3Ndg/tAL+NzGVk9rYRuGB/Um2Qxz3y5DIrW3cEDnUAQl+JIV0oH7uSrMv0uRgtW
6+LWvqn751cMYes8t+yRO9GYzckpYoKYaBUQEfsXiAJowyIcQ8x4RIJIheqxeqny2LbGKwO+dmzI
5mnL0wW7d8LeC++rfufKaJvNyM5HZULhJ0A5UDeZmqW5VfNXeLxRZh8WItIKNCQpRsDiEorR1jxX
K5exF42EG4uOjcK76cWUNE4D/u7AwNWyjSwVbHbNctDDrVRzH2G+JkFzoWQCco3oD0vT6j79bWMp
uidMzBoKQeuvXPOXBSoTGYiyh2yyp9sSMryGysvN2t01zxuWh3EtwQCS17B60ga+ACTMLJbNFYAY
g7dhOO8PDTXHJzn4NjdKaR+hFUdqGM13ymK0eeEo7zj/g/Mje9xQZV38sv8cC92PhZUGtM+w/LMa
ZR8K9v6i+B8fS36KHQg3ykL/iswR/YL8l7me1onkK+kay5aCJ/cLW3qw26UEdRbtro2r9aX5OnKj
Y2Y0+dmPtOlZbVs48L7WZRWmE06jTxq51J0heJ/gLG8arFM6LyjVJiL0CpLglAgz8gSGj0beL85J
1Y7coN8CYl4TVD50YkSRnAW8U+lmj+oOsQQHwPU3/jcqsYN372hRe3YGl9RqH3xNsI0nBonghVye
BzKK6BcVdQeN6duyNw1BmWjb5K83Du3O2Fv0t3eLNJOXnvJsN4HPMO5Jgc3SH4uyvOovUA4vtsvd
+8RKhDN3Ec4qRYrLPCtSKm6Kqfqd5TXYyb5s35qUkRoxgtBF2I1abGFi+B9mqVe6Pv0ny3pwaTqE
vkAbFwd61gIquBROcdlWUUxDGAWGrObc42UHRlaLnlZdRtif8w8HNmO4vuUawRY6e+uHN5ep1gw/
Z9FhCIud438nbtqztJFlwRKokJd0OJPlGTRYuayJnaXtjTA52nd+ozip4MhJ5GZZDyczXYGdOuHc
HasCoT8qmSJ4C+0a5d2IG4YM4/3sglQ6R5Cx89uU7ahnjn3Xssj2oiFcIaUyjIGZ18eGFlgcqlPJ
aSBfp1R3IUSNEpEr8ECnVrQlivo0B5SqJ60fyUTAoShIJzzNIWKNYDSkpQtEmWmdCmjj/Vgg4TO2
I/wPW0XM2dQch7cNmwIoXubFA5+9mLFRJbyOkJCDE+zncIHp/rj0pUdpYdhOWbD5OJSpVGmH7/tz
00qxHNwh7Ve/+EvAAD+WggoG+pMMGA7Ai1c3miJiQJ7ZTOoR1u8oXOJjaq914OBXGGcq5kTk9AuJ
nJ5Fa1Bzhg+N3fGX45i0sjAVBs28lKOKaQpUa1B/zOg/YOI9rqJvTFUqjtSYi/LrsM/LU7D6yqCH
GVanANfe2avG8VIJY5x6CU4itzwI+Ldhv8SPFkMMDnVTbzVM7Iqtpga3XFden2/56P08a/Yh5py5
mIp8m9z30vyVyGwZz+J/1VHHg1a+4if2JU3i+ea+ebUoQHfwq9KGPKGQe7tK+nCbFbYdSn3/1Bh5
emr6cApjplJcpwYfFWhcMMlOwbBuXIGO0ZAOd+/abo2tACoE/qI9w9gIJmWQ3HLMiZrj9sP4Es4j
z190IZ3iGvAEt2qGX9h/5u9TB+5EF+CIe2Q939s/yOUZcNeszROU95ZE7Oz/g7+PEROlml9T5LzT
oeDV+fNGPFc9qKEsvzmvMfoR24/niia12YOcAC6IQ6Km799cPOb4RATqKqcthNe00nYHiNyxLx3G
fP48OGuSwx5QLZhLwoLUSwvE2MDzJ8PfGS/L5PESv/CETrBEw26/+97Umau86aiXDtWj4we6XhG1
U8qoWhWN15NP0EFosZR7BHqu72IKDdNqEqXm7qi3AFg3+BlaFb9RZ5aJrw3/Gn5lzL+81xWXKmp3
SMZp31X+bqcY+IStiKAXsQ1Dfhi1/eIa9AJI4WizSl65tNvHLLwmYjYjqw3tpf3gTzQuqg7XnUii
F8CWW4jrysxGUUqnV0gb38Q2H0UF4TAhQMLXURocM1Gy+nZGNAY69tTItFNjX6L3J59qmKkTmyKa
6BKmo7/H9D6PfMGkb6BGSI7IT9r8JlUM6keTbunwsDrDPJq1E0uHpvU6+IaZbzHONxwzcEeuz+3i
ezZAvJ2Mjq/vbi4lD3p7X5eJeiNm/ZSoRA8eYOLrdUk0lBqMk7SIQNosij7pjf8B5Sx/+/uyKixn
iCO0xAJtxM5q2HnM+UJh1LO9Bc1fMZuQFLRe+0tKWz+DPUc4rWkhcOKKfq/uEZWX02D2XGRoTru/
g00Tkvc5Sl/PqbuVlu/W9y0L+CgVW+QkAVFtA7Ig5zt16VzjEMhXjoEiOm1Jotwnv68IbezsyVAi
HwcfX436phwj/SncG7wSst4MhddjAQpxsAyPWu2wvrFqqu7V2H4jhBVpD/hmARCnjU4mF4QPgdNn
WbkwaZcXEUBKLpSCQ8sIlRh7rHYjrt40ylxyKhUEri9jYUbrkIk5j4tDY74zLP4k72dIYWC5qrkP
6+SYjH2YDV+YyktZdAjE7m5cGOwXfSH109/7wIjdJ4BQCspb6UwlTdl8GwyzyjF6GKk2GMICsl07
d4ArnMGAe9glce7Vqi1/q454y7/yaSFFAlqHxVnkGS/Hnx53o0QSqVV9cPFEC0GHfeXM+MOwjC5G
Zy9iZ+hlPd7NycOD9/uSiC8eOdh9F0iaYWnmmWJ2WFCntbGkkTAOeo+Om9/AYvIAqmKQCadb4UlH
r0NQSPaxpIga1ZnQpXXFh7JOQ9EtFx+iX/EJ2odEde7rFcHk6u1YM+1oGBLdkIDHIYzhRjVizUaW
TiNIqw6ps3hLCjJc0Ba7LYk5jTUFTKa7ee68eQ4EAMnn88j5IR+3ODWsGVJiS6pmXh0+rbfxC/Wu
c6stYlH+LiKBTca5hlrgBlE+78y/F8H/VMQse3h7/aNHX0liU3Wr7N8GuWP7PBZn9LzwjROng+Sm
0fhrpPTlJx+g3+IKTz/MMmeVD8w5YP0F4lZx3VLrZNzocOjQ1q/QuG975QTMKJJDn9lWWq5oBpVZ
5uLsRcf2vnfFyoHx+JmY27i1iUfD7BbeFlYp3ifbNrGPwzEEvTR/QfpJHlHP9oSzygtmXdxseNHW
tSbCCYromaKY6bp5jTsa6XlmxqKwofWKHB6thvG0HbdZPJaqKBaXdFYzINzFQCnvYpW6NH3AEEyL
EkiScqbvULPc+kZESRqefDl/K0VErZ7uHMyE3c7UPDPl5eyo+1QZgdbdsEYbBsVkdPLKqnIip4RQ
GxYPWcSf+aXFaS+epWyHXn2fuWWP9dMPa+DXKJ6Xny23w/okDeuAHZ/t2GbRcSHIYWEbqJBjnPnS
HnTSVs2rYJAhgs/tZgg/BNDoPl4ugnIXiQZW3DKYg24IN9FHk/z2ajKZ0yhhmGeYZ14qkaozlwvO
Lr0B/67t+R/USfBlmOIT3qGwKKbwnsN1s/avRcIfzj9/MBIjbRjKFCpd7qzZ3g0U+O9s31R4u+vQ
rJT6nqBPL8ugCGgNud9myyzhn7NsZCZcYSDh/Sa4BFIxg9jiAkgF778CgjYhkO9s7nZJjcIw4RRX
pslwX/S4bcc5c986tX1VzUcD2E5Dfz6oq7aMZFHc7xle/wfHPHySVfCFqdwj0G/tRYblNKPSQznP
66BOx0vHnQs3rCOSHS+uMCRtXPdnd+c3Sxxrt6BDNGOSCEB5B/Ta2jLKc25uEks0lgQb0nfr4bMu
AZhV0YXmvH1b2ka46YJrkMvIDtymmGPAsuIxchAZpsLam+VB7j+kFVfxPwQpgoRCbGtkPS0LCQR7
4MWRpsgKyHaB4kJflHW7GmN9N1snAniLvtzO88iBnYJZJGqNGe5fZfIbTI65qYkO7mK1QWYZKMYl
ZZF62LW3jshgkKeYROAaXtLA2UeBZnT0FQHMQcsPmU2x+VWCatlVhkMrFz2rFhGmb0Qm4AQ0DStI
qhKJYahct8ttxp/1VIuLallX52/DmbtczoSRv4BHbjMe6c5LU0JnnlGnY2NJuzriXTzeCangzqzH
ROu6V6abVQj3kzJr073EU73UTkwo6rjUtDvqYs141vkyZyahQv4Upjm7s8izZBkm+4vP0j/ll1U6
l3WGtfH6Up2RAn+ZamXzxLQoPuMgBPxGyWgtDnR2PDobv7m9ngreq/sV10Vy+RuL1mVsGrchhTRB
GOfBkoHhfB4FL/rQ+SFUVy3a0KACC6JFHK6KO+Pte1hndbPZ1ASUsnSi2HPIVxJzHeuuFS6/ld0A
69HCZ4x04ETdQH/3sCPHhM4AJfqAhT2fwOgS9WP4sKI3+FQmHd4hDVvgeJ45WfbPEp+WD6wQnvLM
gK3cbBB7FjdO2BaW6KpTDJBLV74z4Qu/3DetrPxrDIkINpyb9gRumgTDxR5okFTmGVBRcbLoNeBQ
W6gLoPGy86ZHxV7J3JQuA11KX4f9Vo6HPQsv0EYJCvGIQ2qnC5I20w3pWuhVT6aslXYLltM5bR2Y
SD9/VDeZ53BtNOM6osMCrr5Vd8WFx1nlgxcUyeFSLRX+LJ2U9XDGXhfDa/A7xOkf+WQSXtmFc8CW
m9GYl0V7hyHe3PaSMdbUTbGWTvMzzFgmzIojT5hcI20PbP3rjvnuHnUZ4SBrolZQxPZjyoOJ8nSE
pmXBDZRxddzQZR4Li6YN3jkQtlNcvnaW44AWKs4EazABFXfzaOCf3FE9wAJ7DcR52bG8DgqfAJV8
sV1ahpv7z3BmsAedJ1ruAwoL3v+nGvhtJLYl1sRFyKbh7T7k+20KhQK5RSdey1VsEf3ZO0aksgbV
QF8M7OyLJ0eGhRm9d2QUJH1TWZ2yH7FVVXiXbGhiHyWkzN0BiXGuEXQyfG0pJgFs6LefjlcqErS5
jqyMD04wmX0XkaIkjlWvMwV78pQcUf/1zMbngomLcKHVcfsTXsOT3XXF2Y0ajUUvBKO5VC7GhxBI
QTWDdkJAycNrS5gowosbmbj3Lgz7QXPWwI1+Mi+fUy+fmrG0nI9urPFu0FkEVvWI5RBHd0Fi8rNT
r9nI2i9mcEPGw10M/IVyEn960RqoTrUrklNrIsxqsrmdEaWmE6KutF+AL+Qz8TctUiHI6IoGE4He
Y1khqkmSQRz5a4XOl+7tjFWgR27TkIXl4hRajHk6rugb41JVJdUVrzaXwQP2UlxYFFbtjQsP6HAo
zPTnDx+OtgSPRC1VprHWqvjPPnN9M+RWmaqG8L3fFK4+jL8Lcl2PPSxanu0fP9mu85q/EsaM6hGY
MQTW22gdxEhGwonXPBV2mmyqYAeKt1EXrdrFf8NW/N3MPQkT0LhdJY24bMduqDqrd4JXMlbCWly/
knkfbiFdfHE9L46Hc5rTKjUfmHPeucu5y8MYSmsNBuHUb1JEdiiCWLz1DJbA4hrX/t+RRazj52KX
pWfgw9Rv+pgyrMiJm07dlV6yrG1JmVuBuQmCYtaEXbHz4rDRXSiYUCZKfOHZ81xQnlApOxMpAELP
pXJpm+gJ7Yb8TG9nJR01B+oUArJbBqQFFhOtLZABYYxqmK5nHH4nullABxwFtTMLGJX1OLgCgyY2
iOM9QkzVHyJ60gSlmiDPme2O6s1tgIQs0kegrs3XVU+9JysjXkaDxlUACAghVwj+AUYrX92U40Uk
t4La6MzvVqtzfQV0ICxtjm6+dVvUNg2zbMzl1ExuFFED1pXLl8kO+l/xIsnMlasaK1B9So08YqBG
+S4eHelY1Z8/ve2SIlQKJRoHPHdzdqqip6nWxTcodFGaXSAmnS0rZwvtr3QvHhkB2raky5t6xgV3
eE2VhBLo6aC/vPJxtmUSVSIrP/b84ANUF4Q67k0moWQLs1aFe/jRO7XCkc0Bl1W7YVKhLWU+F/58
D9HbMXb5I/GsmFsXQb05pPjD8VempJBk+7whYO5xYskVJAVF5kGcOJdcoy4M1Y61XoE/0wG/Gihu
I/7DRvd5BFRh7Kv/dP6IiwNGC8rCGlQWW6dsvZVGxeZ8I/UdFc7nbX2gs9w64dwtIa4xbToI03Aw
es+4CpnRErxyNu9BRnA08sGMLC74QBi/ekZ1FXqUHImzzvvAz0r56kHydGS6vXIAn+cK+I6kt0cM
IkotXlbVA3r5nQ8pQn5FKTO5WESgsiaT1OTOvYaur8TILCXr7ITLDJmsaMoHre1OyxLxuAXlNmvl
z/ytFaLCQSS8AmzZURaxdne4HIeQJaMnM12kOHZYgmzMpcok1CdbT6l489BhCZsoB1ahnKuCvqLT
YtOU7yoi41/Xo9cfeI+Rzf02O39Vun+xnVdcSNl39AUaznkTFDqD5Obk3OchUxnqvKgK88pjnL3e
BKyHtkKjEsoSCcdY8qjGZ1InHcdleNAhcJc5HiY77D/l7B40Skup8m8V2leX8kLXdL3f/U0ow+/q
/b7nkwOV0B36ylatJStdQbJbyw7YGoiY5ifqguF+JIB8W9L59G6mqgDDzvGk+opXwJhyhJ4WZdjL
B2iFGkGoslANiSrG9SmG3ON5RphwO26hl/7HaanmsoEWzRlFA1+nGQ+cg0P/LOR2IPEeJjp/O/iY
7l5+KmtyYTI0u631sHUfSYljae/DwLCJRRVC2wJ8OdCCnG1AyCPvgYwjbfc+XscgPKLDoNZuG/0i
+Vl5r8j21JQjjSFFxv/p0Kr6QUPCQU8FfvxC03MauVsbtLTNmCp0imCEkJeuKw+uUUjmx3cPEdjJ
8i96nUGaHfZOpmepajZ8gI8lM65yOI9X244v0aKgL8Xg5EiGQ43iJrC+6Lkav4rmKYw6x36wfWXu
+zgpPnDbfvm8XN3xl1t3Ws1H54iG29iznrp+AiK1wm+NIUrcM0SErJWAGQALEyGpbbSh9IAS57Si
s/ge2jDSVDTCKw9z5jTfVR+FsF/dZ7i3mLkpBAIEEwrTx2TGKVp9RPq/WD3ZpF+TT1D6PDze1gDC
Xh+kqX1lWOWonXxU8namMnxRMsbHs9PP/fdbxCNLj5BjAJbQmIsjZEy+fa+IQCgfOP5YjDc2aYlg
RAH0MhUfYXE9d4e6HTUfPVYgAN4wBo71B/H8qBEgRs8m5igJJjabWP1Nb7nKg0HGPXPb5aaTnpXf
yxYMjrr87w+MbKQyjjn0Z9BiJoadwGixX5/XJb669wJkXcIif+HipnWK61TyW5V5uRY+38hpNNtR
Pd0cikr7bDVFklo1RqpJ5xLfdiQE0bQnmc91hpVgrnFj9yqx6xPVR+J/Jp0DjjDMOkpiFKmS9gt9
XWdxYFk+WYPx3Yy4TKzqFkgchXZQpzFZJPbreEjqpuisoZqoIjnLVFiyOstvzsrbTVW8xCMBGqhR
qRZ3mkCHdALXHZ4fBfRAgl2nFxfq0u+x0Sw7PCcxEI6zQ0ctQALYsVgpxpcrT1Cjmi4kdAVklUG2
sHzPvWsIBPfnVzqFZVVg6Tl7JWE9CHRcrrECMOF+2Am7yUyNsOeSrj4Z7vkhZTLdEJaiuggj9VD+
l3YU8vE0jOJKFJdpXgkZyNqTt+wE/LzuUGJcQc6Sh6NLNeY7j8nPWcoqY1DcQPNGBr7OS2TRBYgY
TGDwITskzNwlOLE0cI2bewuRhjbllJVJytBg4eJTxufRMikZsxGEi+S4ATtKW5XTynhINHeEwl1k
HJCaO8D1dLMm6iorQr+v+waU71i1wsS742kCI0Lj2Dn5Mfj3f1j2UE2FQvcCQ0Xw8eBeyyx5yufp
I5/A4ZoDt8oWRcnnX3m4m+umOUxq+j2rAvIXlg17e8aRL6UsPR8oyyx5X3bcJ3M5HWdZXe7ZmR3t
ndLxT36IP308vz4zEjjbhD7wShbkJwUx/SoMQr17plnHZPk12Dd3d67VfJy0hHHgSc7tv7brUYKV
rdriYUSC4f7fszQd0fyGygy5VzlN9cIEVs0rsIe5MEjw6yiNqQYlNQZHc8PL6VoNI5ATXIsXcEys
GcPjGWHkaWRNIDEpEnaynnQispDLGFkOi9clyWwxb0BaJbRE304EBxnCcZ6n/NaxiFjGRz4DUCYp
M32JT1Q9kl5Bve54jVIdnmQ6E6E2gCXCY8spmKBnTbPqofbtB2ArTSknr2lpcqEYrBQC31FUwfAW
zMwTwwggVq46kETXr5r802tQvrKMM/1QX7CyngY6tKTHG1wGiqGbi9prU1S0pzPpxUMSi+ux3BhB
eptb9eeRvnL7+nRWPfjMpu7aT1p5hNDEcFSvxooxo8uj2c+l36bpSY2U874oueJyWNT6QpaHrnO0
8ub4phKdyq4YcxZ6Oye2xXdBzSWliuDWqZQpe9qMxTpGvPstOJrKOxlOz+MXAWlVwlgBPdiAb7w3
CJqh1A5ErG2UyA/Kd80Mlc2+YwPqQ48/LZWPpiWZSSU7RucktoxsUqwyNVfG+HRxEVmLsGayxYv6
1HOF308116y4ancbbFrOczZAJJP9dtcamOZTFhzDP8npON692+DaYCsWQ1LpMjdFgdtOp/HdlLOD
c3pSYTpb9jqR/LUnA5QHFy6F5/wJt+7jKGWpA/DhX3/msrwRYRJPrnjFG7OX8939DNPptvUulp/S
UYoa8Szl03+EWFqAXo/QzRm5nc5li7GRPBxa0+VxGZuj23hFXJzkQVKGkz7zXjmXniB6g4tzR00l
oNb5I4MFpPIzIQGotcbQWAlr/x4vtmHlEUZgQ3nzB0eRt+lhj75Yvgy5c2A9EChlJE5rdI1g5adf
WKoM09seVuvQy6cd0FqlSttacF9/tEiCo/HY9PPO1gFMTAX/NbvEWMmObjrno0XK2WKTR9GCkeYN
yD/OdQjINKyB3cpspFHiPQt1ABgitJaDf0qbFg7qbeaCPk/oFqfuvLLbLfnavrJrZm3d8KAzNkwT
UxhK5B4rVCvyFlErqU1grbEfQzeJJr+i4lcIYwmK1jZhdRL65UUeXsJRhnxRceY7FdXnMrNDT+Ag
M9MpQbDUsUe+EnETqVVwbYpTWgy7Sl7GmrErj2Y/yLNzsaI4aQgGaorNinw0V7VfLaHoygRMIkfP
El2RGvZJ3wkrUxYP2Aj0ZBM9XVENuAJFb7MPhXM4Wr8xc6shX+IVrTmRgpPBwMzCaXht4qTYozNb
ounJObGtLmcUDinZWzfnuENY2iiF1/5ipq7lcXeOjI4TeB7eg1PEGt6xfugnegEPZ46Ql70c6mYW
Ub9+281ewWK6iwmXvNrBb5yQACBOz3CL/qEL7tRBNQW7zuNW095lrV0dQXqmU6/Fx0cN1RBFXi2a
ISwwdfVr1c9qbUmtt/azWMWIdIEs+sBCcFk4+2LP8g1EtiYYsKS+tnEllBHPm2/spedOpeq/m1DJ
AqYpAqiNCFhB+2TYRf1MnOH3a7m7xkfBy1Jt6dC7zNARKIFPDDnt4fW+LSK4UKujG+xLMhoQHXWB
jKX9+ND3tTwLOPC70odznGm7wBy+ehWMZ0BBmFfm8GJ+I4zPn71/kwJt9zvq39bIGZnUJbTNdGJV
JMc6eWLRXYUjr8sl5/AU6OFYJ+fZj9fjHafEy0Sj4w5J9MNuNeF0+tdyMFdjS4z7gKOyhhMaZvsD
WxufLJF9W80xMyqCL8nkvu+Bfs4Pq3BldedGB4qIuQBJMUvJObg6eBxChTduria8wzsns4C/zphJ
UB7gQ1aexUC04QY/4EQv/qMUJDaMZS3rIpRnwYWbpr6XbRFttH2SMJHj2hoYIaqAoveGamomFHfH
NsdwSOMIGOGUoiGmEKjFOIh58z3i4SyeRarPOLdrF3G11JLsr8whIYjCeEtchc8TYFj6i2esRDsJ
rleJwtw5ewLC++oBBREsAtsQgyq0dCEB/+II8eeWVYR4LhOb86636xo+Xs1ImVr120LOmWUiyhjy
Gvt1dQF5OWgZZEAa/V3oKgzP1iE2uV54YR34MAB12El+gECmiFHJQyu+3la1Eh6Nro9bdNSYpSb5
Q56rx1vC26FLcbCQZmNssM99jSY3av25sEN+Kw6F7QPMCcngm+4pALNl0dkT5he7kiKbSZuEWYd8
IfCx2pLJAOx6mSATj2Lu5L9Low4SkQrrwM6YYfOqPnjTo4yuF7V6EwKrDUyjDV8m2h2LsjoWuavn
jPTyBeeiT7jmbmoKfObHUb/sGE3pFFVYIpy0wgKAoOLt0f5Iy2JBzhGiJGs0Nra4sq/X9SiGBwPl
eZSkX+kVdR/zdrEIqlM0ZKl+257fFLJDnIBQ+Nuz3ZNP/jYWoflIHUvdyl0Y6byiwbD2hHUYYUW6
cgzRwdkcMRX3pa7a+TAO3F7Svh30nkfgW+SuxPHcHSRzSfnQwZYQefkNGL13SAkek/NjwKvmXkHx
NIoIMQmyL/CmsS2d+mk8K636kmqCGx5LEEoADlwqDH/uFf3KMWap9TXK/fqGKZ/dFvWuMUlWAdAz
0bVuvIxR0sGV7NB8tKm4CmrAyLJRyPgc0jkbzZU0JERAnzIkrL2wvkK/kP3WtWzf+ROC8pyrgaTy
9A85pNHIk97BnmQn/nAwRbio2G74dhExQdOasCMaqeHNj85+RaPcl3r23oqaf0udiuKD+aZswYd3
a2413lVbrzhU3lVHe506aYfjcnvW/ekZLYB3/47gzANHvl8qBAEB1Z2nhy0rDhMPWqSaeS6A7jc7
MfiSkBcz4B2jZunlMLUjDSfAiQbIC5yZW3ArRHyhKrs3QJw4bsobXxwOd8lQo4VYD8ttxpigcmgx
jiR0r5PoSQENfueUvfps83VO3HmSoAZQP1xXbEcnG4kM+kflsoFSRsZmwa/BusLmCHmSgBE11fZC
SbunLC2NhG2Pz+GNy+fkOUjjgisXNrlvJTz5VK0Gf7fUemrQgwgrEVUGE2j/Nf/++CSBVlAbCzTL
/pgr5/E9K2KVOlStYIqKC09RuLloFLiu1gxK+EfIGu9SM4kDGB+QDRcU3svY3oz3203X+vK3fQJm
Z7wblMGLgo7oeiPG1s7axLsFJGZGqcY/IV5alFozjkuf4mym+dpgzNCTXupR75W7FY+vhNKyrWgF
8poEyU1DDbfZl7mVb9cUrcYuIZzMmcQLknSTGBx3LL+6d2FJM2+YMw6N7smHnNy+4ChZlzKPtVVq
sKYs1xji/2JzYaWvAqTTSrn7mXQcpXicXpLKxGpAbBf8ZvzIuMaoAOiTfFmCyU2fsirDZLE2388N
Z0vG33ByYSr154i1rsy/s2migyTWs6xLSTfp7u5g48kt9/JwUudfMSzgBD5n50PWoOJ0MuNrM/vi
e39hxxjqg5osdQKWiSWt+T2sn6CXuHJzK7y0bb3Oz+5Ks6lGWlVQGFZMflsyUk7Ux4KUEyF+EW1Y
cOGVIfUc+TLVxatTlvR7IT/hs1bHwR4lpAVOtMa1WSuFAhbf2Rwq1Iuyo+yn3rGr35uxabXuKCca
7LyA9NqjZW6zaOoY/JkO958FcJ1p8DGY+Ir1AkKHCQY4VJW6H9eezWupN9OOP//Nl0uUbQ3wwG5V
7ufZJV7xQRzx6q7BeBoc4PuZ6FY1OHtRwDlMnsziE5u295CG1j7meELxZX9NjY0P+Ofyr0g9mvyH
IzVjnTX0fwZIltZxJN7fTL0E8ekdhp7U5/TcYxEjOdgxZjKVd6s8AhENC+I3c1QPCWUeo9kZvinu
xvJQiJih2yHql0QKf3Y9ChX+lVcJjl7a4f6A6uTdyfXw88DMqb3p8sX2Bgqgum/RRmyfeNK5h3IV
bg1W+heBXr4YHQqV4yNPu3zfB66PplBzKHGWHPh+dO6vb7g/Vhq/KGewATfUWJkWu7h31flBCywO
96Qx1GJEhqyMXHcTeBD4by69y4WdpMvykSVeaGl6jBGDQ+Ft5aUtOcADREiHpzYDAzOmItwYK/OC
zCOwRks0TQ9cpl2ZZ08RnIHbXs+En5gbGNoTFqZl/Ak0rV149fSHYvvpupoAb3m10cZPO/cdFkov
Vmeixku4KMC3XsB/LgjOyHBsVbRrX44D4KD0QGnOkjUmGMZByyBLt/X/yOBvtpM+4FmJntNRTcKL
t3rSeqLcgc4ObzFoDX5CvQob49Q9mypIGsGsIbCHFIkzAv8eMZQInp9dOrKrwN4lj5eISPjUUHUO
82sdZNmNkgzBJZbX97MfYHHqDGPy3p93de4q1zf1N8oJoXJNA7I5L+z+ULvmozT7/F15uJmEjJO1
DYyw6bley6sS7bN9an8PHj7W45skeVGUPyeEHjh2H2+sgm9xoLn1JZNUNW3lOjPxNtC7uWEM0aZA
ukVNY17hA6g8vAawGaZ2vJ/5po+YGbS3zfxb8MluIdVHptmbTNN5hlB8xAPYliuM0Oud+qhrjKXG
rxWEECfyHY2x1uchkbSr/xokP+LojQp1bjmtlnroIQF/SsP5j1OYHEfYrPcSzoq5SwLs0wGPrOcc
+0dqEJpynxOVY2BuiNd2hIjt989uwoj5eSj0B1vPF3Ou5IFhzEhlNuPPbVQV8WjF6suhC1cB/hEu
GvBSeLBzlOr6MbHxX1iJmPPnvxjm1gGY8HipGstqBuGH0nzThcXgVKpuN5uWiPap2RGBT2ttwc/0
pHPFfgw6i5A17f1g3QKchDMgnVFONUe7GQYoWDjPvk49Fqndn5riTumhL6vx3ngZKU7T6TQGdgbq
BfM/nToti9htrviAUKp3PN8h4Z7owYX2NOETFK5lb15nr4KZRJ+6NbDJd0zA0zs5ap+bxGmSkSF3
bP0u068RRNB+KaiE/MXf3xOsX/BQ2557OAYaKEoEWFiEYMl3kkJi4Jk31+xlCFKy7qH46n60hnef
Z0RPBoZCUY2enW8QrrftZNwCIJ7FRz0fGsMdnKnCkYinNbmaFD2fVpebQUB5Tgx5DgsOesxt9+pQ
KwHXw6L2ZOw5K6FZf+dFphgIZSF/IWD+6ZAMsXoNDjgviIQMsReKPgt0qzr/6Oz3v4JjxpxLQ8My
P2/8T+vxnTuo1dyGeNLBGLTXbH85KWbjSek4tIthzFGzCkQ6pLyU6hKINzR/q8DJGomu05SOUWIp
Q1LKbt28iYDAmOuOrnocV/Ad+zLuTC9pqvNjdB8V+V7cRucXrvfMHB2nLbQgAa4Buhdv3r/DwIO5
0wfCGsVI0/1RwHFyZB0hmqNK8x1JCr46XGj5HKGBvhmv6kc16M860rviCbmqFBBxXwZON/VUaCfE
f7rSyJf/psiHV0RXYS8KLqhFItPFNAanToGiMFKD/frbyQz85v9T/wxFsvrPnaFtJKrctjfp84SH
M2zKuHXskP13DBGPXrkcoUI/2abykFg6DqMAPid/aHRW2amsicljIVQmDm0dFdNeMo5ZNDV9yZuA
1EaFsM+m5REC7N1TnUSDpcbI+qqWxCxsh+qp/TmWNgQD1OevMQ6U7g5PEE7kUvI7dL5FCdlhI+lN
dctuGaWW4uyyBmjNYPhefffv6cHh0T7l6VGcjvHazandKB2HeZsgsjEN0dPaXRgWX2+JjUVSi1FW
Y/5hBMCBMgAY6hSov0QGBup0doVZWuJM4iEtzq89sufMr9jKd8Kvcf1oZYzyAu8mEO7zrY3hB1qt
IlV5edIJbIuml5LO6Q+maMpDtpWF3DOnMV4maeOVZ7AorKtXZKrd0a3o0fc74u/J5VkTpMFVWzhZ
7ivpK0ZFaCbTNERd1TbdYB14zsmZ7gWP7voaaBc0gJZRUEsgFaMamqkEP98pr6l/TmBp9UUi8SjL
SjMfypMLWaSkwAFjwLEjBeMT8vckzsW1obduDKRkSW6l82roTfRZfJupSpCn8/DF7cXxIkiS1n5t
4AeeHJwOlqHpym8wOXHWxKQ9cypDOMANVKNyr7KHViUwDRwvc5pf4cIJcrwSb5CMTz9cmEbF5JFt
13r2PwieO3eisspQIgfd9dpigWL4lHNMtmQKRpeQs353Dwu369+TET3dheCuJ5qa+GiQV9UHryGD
/mPDNjt4Kh+s7SF725xhWP8ANG73Z5tJHcv83sKc6OtrPtWGHa0FEsyDzdaUtZ1Vhq1zVSLiioA+
Fcyln/bw01hNxl7ETQMx/jJJiTMPCtG3j8sDrBksQ43OExnLC0PCpjhR7DRUxTBZcwi8nAQsTIUu
fYDeEBYkjCLik6P/BtcGpvEOReZdGDavlxmlal6EQydrpjqXnUUgv8SO8hshtHgJELMqC1Y9s6IR
aO866f7oRt6NMR8l7cUhhP5PvcOUEPvaOAnVou1oK2dOTX6Mq9NPf0xKXClnrCkekVBJ1MJi9ERj
/3DxZxJxWbYRqm2rxoYh9H2lrL3FmpBhEJq+7oZOF0KSXTfgcqAmvNKW91C8qxAMSJHjd/4tR9Kz
cjM1n2DO/rVWmI/1+RlyGOaUqeHPVd8AncwGHjWOmC8PaQQKZgtvBbaTveHzXRrgbS/MGtZkPHNa
VgYeVr8BLdLlrGAMQGj87Lv+bujlpVYLVpPb0XbWNwjmFqbK3XSn6a9nJ+zUcj/GY4yqTo7hqlfg
b6pGRFJ4/8im/36dgBt0CMJrzFNewtd9JYhitDcgw1PlXzwm+b5vC8wbEy9Lx+TXLlf7z8zMP3JS
SkUp09Rwjb8Fh9cuKYT/468CAACrLrLtOevKUfu3+B3VqXhRjnvwucQSDgZcPvvB2OdNgDLvQWGi
m4TUhwUNbGd4qwzzgvP1B+G62AtW/oyBEVf2rReuSuW44TEviqhPdDzSf4UlPlCgNaqx85veeHQp
/bYt9lbJn6Wy06dQIjIdmYnZqx2gJqYMEV+saR8/JctGJb9muCtPrPy2PiXvdwA+/QTjdIfhqmE4
F4znG6/J2pZbDSzpgRan0HT4SR7o0pptIRZdleqPQyuGSmjKgeMRPXBhpW7mZrTq8/B0Vj4CGZJj
f1HjepcODhWiegJbLrn3jLtFf4JkDC6fzppPX8kOrq4qVYu0DMC/Dt8Pf1VdRYOmYvKqNzEMoack
Fwwq37AL5qZ0SZ5nPzFac6p8IEnEqKPypF+jnxpAR+8Vn631Tc2V7/I7DU3kMcQ7rw242DCVM37y
HXO2kgrzP7ltg9UnTiJmDSgsZL2/lOnObpggzjPsZTbA8P4fRy13xBl6QKqawhw9Y8zhwI2VVq6P
DsOyif4JntTKAbOvOWMuRg3O3OQSe3DVTU5qE2jPx5KcgzUxVIvt+XzC8mPyCEtYupJhgsjmTXl1
KVd9TD01E/p/cNdZ+x8w/uTEnABm9uHcEZ8LPjqjcyB4MMu0lysDFQTg+dOBSnKxqAIUEFqRp0Sx
RFCD0Fur8/OF1LEn52FH1vWXF6h3RRQS+18y5dM+0Eq5cSmeGPltIxEU5apqKTmu0N5c3oNjTjT+
9dBIytF/TAdZGoIo+SVRH3dCYznyNdfkRzcuPADE2o34+lksaZeXxcAmf8znfbvM1R0E0na+xYDE
V9hbJICkcz0Q63DQVNxlVdUhk8C2KrqV3MmFED2aLFPIxHYmVXFvA+96TaWmr5FVVKP6g9zqoIqx
WFp9lrxiJOOKKRp9glkall9W9wn3vYzk5wty/y/H+dLfG5py+ITPcmvkVpzJ/v1izf5Vp63sVd4W
bjJU0JctMmgnP9oZVEUU8WWTq7P3I5t3yRtzwlw1dsLFteGIdP9EqxfKDCpxsIDIZQn2M+iGkiXT
XrOx4MAfsCC6eEHU6zdWlU8kRyUFzBgwuUHu/lfGAcbLbvnDv9rdoAF/YHadmS4EfBx/Iejl49UN
TC6GDDvgqfjdSuSv2+sNSyKEQJ5RfvQPau0f15Nw/bV7bZEXPHpsqKZZMqjX4zgXpEURybKst0s/
M+mLvQObjXt4q06wyHt+Go8eE8xYDeKZCG+wEqXeJKoS+RuniKbr5d2zEocd+9P8tsFCGu2xvBNL
klCSumJT3hTRnZKVXxVoGDUj0Wv1JWOC4zOXDNG8Ki2X2fU8t5LiQ4Vlc2T+c+dEihwimQnBAx9h
PQtqExcMVVO6WC/V5wOIfOd1BAham2QHPuvHjaMvxeTQnRAx8S4zSeQ6GoAg1O48NMUdZw0MCa62
0ViTjRktrDwcW+H8td0dZEyR2xfqrwWpdgDICDxvw4eaZLqMHYfFYFr5U1eRaCfq9CQwd4NcP5sB
53hhC3loVIDqLs5ZVT3rEMYJjUzFYl7NU9jQ84NTt41FFwfvXnFjO9WMnS2lgbxkjHCj29ZLaZNK
ogFxygoqiiUKjSRTd+k4PZKTooe31pke3G5p0Ss6EVQhD36ELqMefzUFhGRd14NFtpK7Ow0dYwDJ
07knj5LQvVgI3ceDQgi6fSTA6yydJ1fku7y0L/K57rRwFNU20FbzeVtkZebHS2l7EybG2Fnddb0Y
UvkKU8/jwngAg2reC/zCG6Xf2FrSG+xiW0HFFRdk/ez5qIiiAitzoWe6BDYHK4vyT1mL5mWB0UVL
gbfBoLpwo3VjzG7ggYuaxBsEhF5jITDW1xrNQNdoZgrB5RulPg1QTnfsgKrtIZZvii/j2lChMX2S
HuMGdG9ZwqKiLIFXz4lySqd/iS1G1BZwx63z8fZcRj7+fciddfU/YTnnrx5+w13yuBc5ZkUVjfo1
0p8XnEafkE6p1JVc0VH9VTW0SUlLGhK79PLfTHJqqH2FqmGXuElR+22kQvw/MEBwbcy8Zmj5a0Pk
nwVQJ6ykvONvujXMQiCKUO9cc28TPi7gvNVKr9649O3pKFAxwjF26+DKV2nmP4dXphVglE0HAnmW
Uq8Owu1xVO4i8gJ+p3wzaC6AduPZAg18Idu+gNoouoxgIxbaozKsuhLqvJEXNAGGiNacmoBRDcBq
ypkkhDqhcgM0EwJRnoxsfvzBoTEIeC0rY13bkjKTgZaRdUDgvctd34X4tqTIxzqJYqqPx32rI9WW
qajzYqZ1ig/MBpe5ttcQMatRQzvDeL2sVOyA7eZFEKCXU2n8N5043mD97yP9t97PceyLBQbSbKRS
Invl833/sTNHbxdrtyeP8dTOMCVDmuVuTtWlDTpEXQtxbJuGPMg9F8APeX0XCtcghH8Sgyf5JYGK
TPagPVEEElQPGdI50SbZL9rnUBRMpHD39v45/4ge6RyafQGFE5ovMWY2Pzsudms2o8wapQXnxWBu
5vua9yjOFC+EodJzUSKMr3b1WhyNwPqfPV8ziZ2BvDD56gIvnaIgjhzt2UH1boSgLyrGWQtiW7QV
2pjW2lbY5Csm8WrXyRSpWuelC9yvz4qOrw5FGZzDrtaYHoUDC0pPid5oU2OqSHuOOdW8+xtgHz+W
/Ei7hiLOxvO29zJAhOsmjqtsEsAyaXrblZwD4Bo+ysiTCpxoHzIQWO5l59aC8HVZ+s6qub25zn6E
uf89uMpXFRsebzvUUUZB2lZGYwthL8oOFGr1WcValDVzMTuwYxY7Hryuj4wRshHsBXfAWa+vR6XJ
kPDfrVSlMJum30vTXOA0mEyi1l+PJ/eMyLcd0Tevui2d2lYo9pjlmKimfe2TsSp9GtTXKuNL72jf
FmmRW1xdbS2jki8PI/qy7tgPgh7h0uzBw9htn8YnjUvRtQ2PqItwPpBQbt7bCLvQqlrve14fu/gl
bVzBJ1Ndkl09yuKJQtLwwS1ZY4WptgiX+Hnj7IEPeSab0Hp5DV4g5onpditzqE8gUkLOG7cspk56
SxWpusn5yLKh0cUHULS3Djcr4NCbkLLqOtAb39c5PoIDBym31jwGbN/ZS9V7IcfyF294Y4ewT6oj
Kr4OhYELiv9xfRVKElpzgQxhEdaBcor1s+V32erPktafHPN5hhq6W2A/WBuDxPkdcwvcKeeBHVj8
sYG/LwwRraYqJDnvzMmMKf9DVtGqfE0jewoBebYUCAklXVXIb3mBEDDcE2K2d51toZECNq2QizGH
+o4dCSV6aV6SVJUgdO4GZ7kR5ga196dKqDdTAqOL23qnbjKBrjSfvmnQBY/5esWZTtnS/EutjBWi
7ItC6A//5klL3ZCo037+x/nnx3ewnugiIPom7LJ9pvE8iNw9WDIaT/+mAf4yw8gk91SIC8T5QnKW
E4Xr2X+WyuYV9xXvY32yZfq8afKcc7YkIvVgZOQdD0RBJ/5gvm7wpPnHteUv37CpiyM2L4wq+sfM
qmtrEwlkQS/iXcPe99M+F2cKObf+f1P7X6MeNWaIg3lOqy+1wpFAQdIiVlfB1TZkgLdD63Keb5co
Op9QhkQNHTqlBfFJCuyQXC4EV0xxBJMtN+hJY4wNRigil6AqF4RRzxZUPoUo/IifzL48R6fBO34c
MEqoHO7uvLw8ewCHwcx+Tg/c4T4LmTA0ua1a6EZ4DkCDHOvP3EwZUX4zCnV1VvpTxuJyjqABpAyL
n8A92qrGkMX27LLJ1I9W5IJApLbEH1agjDoAA0hRRsRrQjxOU65HQ9lskJeiw8ob+siRtO+hyMmX
FBaZhvIsaCnPwIuaRoQ/aYCzqbDemUaon28rvJujmkqFGwCxPLK7U/mK4ft++cnGsuRCZBH9Pkgj
qNIG3r6RcFXTal/UuT6b+voPRpC35tTvlNYOfwsjE7KoM8gCxBKYr5eWPAIuSNuzGnf4urIr30b5
KWDBJDoR7mZAPyuNQ77NllIV2haw5PCe/GcXHtYb31Xtw573IDC5i7pPf9kWamKA2MpWi0uOYLiV
PEGMFamiRse+BqC3PrBubkUzyIIHBiYTV73zMp1rpcWZFmAeL3uO/offGxSVVYJsQ8bl2vMV4YF8
vtmZPe2EhFZak4y3de9yeRjO4OVE0HPOKjuLTnhcXCixjiaY58dxcVHBj2OJrY6vtCmXbZrrZbk+
MU2LTUK9Q6lp1ls19fYCBACKZORRw9xxyH1x9wtU0nabCe7M4R0sgGix4PzVRUtmJWRBEPcbquif
qP2Tz80fLesVGSL4GPcHSDIfGbItf2Ee4XYS3qQgo4oncjl4l/T3aK/V/9S/W/9q9gaxcWLcmClv
HI1flvX3YNTywnjOJuKMMOC14nYnHQ7vzV6P4R5a9VaA/NjJSeJSkWbU3OXo65x97W9E/x3SKBvf
u7192isXM2uUcfvR6PNHrGWtMcpiFcbARwviZJ/uA5uGada2TeCklqQuY9HrbY8OBzWIJ72sn0Bg
AB6uhbv+YeT2bt81gpAbSy3Oimk7upZ6HDeqQvDQ5KwO8WlXCauQit+ImLYBdXBBJhHTbuWU9nn7
6BdDPIigZllx56n7/0nHAg+U31EtVZPw3q92D4OlzYbU66FfrYVbQzf3qp3cKNohDDVQ16P2G7Iv
VbKCTauVzdDzrkcgQs1fQnws7Wq3Qv7P0BLywjUChazsg8/OJuDlQwOZJI+W9zQpGX9ICqmuj0nS
l06K+xFLPwPlCAH/VzrXQcU93pMCrB2ffZWQ5ygsHWUJjX8O0SnOqfpBAllOA3xFwNKS7354dIwv
m0xgpRPSnNFWWZYR2ED/iW1yKNFSgphjg6n47flJB/HxG6Eaz20XsAbqMF7vDexCN/cg73/kkNxv
LjOkqGKy4t+APHC7km/CW5L/bjxd7YmMu26fztts/nXmPI53vfoQHH9d4DTPRRn/H4aXM7BmZH1a
RjGhWygte19hMTLhEUM7U43xi+1KtcsYrv81X1xvzGD9jEvRvpz9lW6iLTM8m5lc5ot5e0Wmqxs0
YMVL0zmfCLl+C6msCOiH1d9EIlL+GnxQyeXjYT277cJhYyKULJ1ZIbNrVerWX0aDPv/LFF/c6jeL
o4/XzxmxYydE8UFWHJJuUMGuu6mqHI7JIrMzvRxAziZK7BEzGtM4qmQGQm+K9hQIQGX3QNuIQ47z
vn7ICYSexJrbPlnSLY80yGjeNP0bGO3Or6OM7cW2TYtcCRmndJCQDcPlHdyKvXL41eodtkRyNW2V
s9ttZ6I0+9J2M5N5joOSEqHaPYiuP8MzWbkBPKxqhjT7yEEfuJwk26w44hgKa73bkOIqn//K7GWD
5NylDov2GPnu8EpRbEekHpOl7vUvB1C00e2QFgbo6uXvxAweXxZrfz2GE5q/ID+cH2EymNqmBOAF
JTvkTJL9B3v4x0olORn50zWxj9OxrkviOaYLWpUPB3HLPOTZBKyvnb1JXQ/oI5N6Wxo41zqozvrU
8aiCh6ncBxEwkEbexQc4lOmfkYH4UIig2e+ThupcH0V+tV5o/U1zTARLNkQ69Lxbq+cYmdUqXW8Q
L5rBSIdKErTRpCOoGYxco/jdh0U6n9ILclBgfKhaeM6/St8zQsB/V9sHfwSKEW6sgHlUHaor7nYa
EUxKR5NSvxxl/vGiP5umuB240q3Pf0vrvSIBaXEq0TWGuNlxZWrlfwsjo+0D03B5SUjZ3AMxQuVq
1U+qrPRtYvE4kwvu7ylilxUQ27aci7Q84pOqiZF6bQYuP4HfGQUgFbRy0w+3jDNqAvIbdTRFTj9R
2Ila3X6ayJ/3xs0xLNlltrsqjUZXZSh5kz88do4dEJ8vbVy5U1E526rhgvNAUsG55MzSCumhBAzB
zo6xLodXOaTLnW4RIuMAx5CzKlh46MR0IzQqa1f7rLl0f+bsUDEnfK2VLwnUtRKMyXkEezm8sL+Q
eicnHnhjutoyTOzYnlxy6TitZ8IIdXZF83SYq65lM1QyBEsitZykaGK9TXFLcHXL40iMKsOFwErg
s4RogaXLREJjOxMw/q9b/+UY+iuc6BDkrJjsQGotbS4bDVY9Q5brBlLeSOLwVuphAYWEPXdNLQLb
C0oaYG6vgDNPezIidDj6rs2ZvUd3BepSR+KXC8j+KUvWjQPBTdhlhb2Y81O2P/LY6iQn2xaBWB4x
Zj8uLj4Nt/G5UtVSwRbikHA1+FNbnvz/k5MNcEHN2pqU9qD1spGMn/ESBGNSdKv0f/YLz0A45rt9
V5FAwB6LC23MtX0kKLErqKIv0+dvmVVjRnDwqaLGJkkraC0srpEnpphCusUMZH4p4k2rgiwUwRol
3Rd3SmOeJdTjSMHHEQ47xUcuUmMEsgEZkCoOlbGWDZj78Bz9VbiHDO08uAdu7U0oZswFOv6xQw+3
exzbYwFUnoB4JUXDzoVKeE4R/yomPqwdyxXgUNr5Xevqin89dL4CFYMw/9AOXVp3o53Uml2hmd4v
5nmC0mcbqQtFbnX84VPq1GPlTrROk+vNtZ9hSaGXKSOsztqP0SmgHs9W1z/qoPipFEwawtV0J7MC
Aq4Srt2G7r3ijDoLzqGQCHJVAkUaFXkKW45oQoJXQoEamlMwktyLbR+YjJFU7/9a9E1aJ0aU54eD
dyeRyaINEHVB/8i64wHc9wwF2NqLDfufggATJQn3U2TKi6SNjxqmn2C2c3OV5dVZjXLXq67Q0lZ9
vrd63XF23DnOa31L5UHNa2IH3/Skdx1+7n0WU04CAh4hbst4a3XOzDWYvPrRdbDiO+H/wUTNgxWu
RglY2b6wlHq1DaxWyqHYLd9lfKVwRztYAQotmXyFEPnPxQii1TXQ0bf0YrEn98jXv9KFdBvhAoj6
ulIDozeOHVYmYofhMGc0l51UKZt16y5tSaSZwr9ZPw9gdebYsAvWXVrFi+VOLhUS6mCC7NCwVkkh
Q4nFFPK8kdXRedNJt4hSeIlB8BlgRxcWGqi7z2miqXZIjjTtcZy7lVLQi0Fsk7wSL3cEPeCiU9fE
QK80uEvDsSUuaWFZimiRCsfBAXbKC26PvlEyIsRBVNiWvqy6ERVr9yAEjODzuPbnRpJe1ycW71ST
AC3NCPQIoYSSobEf74rDA5iRI7apdq6vTz1xKiYvDCeEj7iiB3aNMRvbah7DUtlsM6JgamauhpxE
p305Fr+waTxUOzIOcYLiYhcv8unmsQy2rajjJ9/0O9wh/DKbABWclon8QX60d1g9mqDbWVjaZii/
FIerEqLNyvkRfhBU2oM7r9jTlpeeIYFLRELJ3auEYLWvpHHAuFjPAqjTSucM8Viq/Gt8ylvs2lN3
pM4QjOvdx/3WsG8zO+bkLM6u+Khb+sfuQdQzfsptaaAQWSkgIGC+Udd/nhZu/fjrNEtqns9SeyO6
zdOUOfmPAAmfqVJWwZ5TVz59svQC04LWMR8DYF6xd1HXuCZYiU93aVVPphYKcWhBsKGSHmSXKcvU
pbfQPzXzrTeuO27kFncCFzVENCzzn0v6zf8TE8Ylyiio/QBDbrnfbg3lNyB9YrYYdnd0q5HSbDOh
6OnjnGI4/0/56iGaE5DYwn91klW1/D3KpAKn5UukaY0f36h/9n/zKcNSy1DB1uvV8JeGrVCcQxXl
vSpX+xuSrHF2bOzurgKTYi9ISiiQWNjeE6b7EoJOB+SWIqWuvIWn96TRvJzcxtKCZw050Zszk5IG
iRaW8kqttDqmswOQhz0xdr7selQAkUqMiNNEJ4aCqKBGCZ3W2y9Gpub3ix5gue+5ACJD14OjydDy
6hPVHDk9E7rjFBjLCYMZkLdZOv91AFcfZWAlMaFI7xBZ8ZrkFiDJDV5LvowinXBoM5npdhtlojFS
Wy4tMqBvDV278AwxcVLHgzIzkzwonpzeTX4YJZeXaONX3tI8OB1pSYwAV/otBN5rzmsH810M9x6S
YtGHyRI8XJD+eKJFy25mxAJL7E4YKmj5dX56+Fh1jIbJmrnn1nyXUSd7M4LLZ8Yuy4Z+18yu5O4g
jfXgyI6TpDN638h6mSyyiLYDrapd7kgeDunsKYrpShC7bmRb3PguXWBbaOBWaLi/oJRVSp+JZyPB
y7xF5sNMy0uDmatADWqaHdqeKdY8eJkDw3o7Lv1CPoGwfrSSG4whCYusOylnnZYfxJJ87vUMhjiP
ED+Kv4uLLBXKRyleXMZ5yhYRY3O52EKo8sEpiu0OWZGEt4Z64JT6lPxwKVtn2V7mMH45Yt8OgOPj
CAOZ33Z4sHHStljeF/iHBzmvsCKH3g+fuBs9hHC4+CkWunlu5/fmTSe2PfZ3VYrIX/pwDtHtGhCz
NTrbIkut7ImrEddtvhs5heOH50Lq7kxl/PSD2M7Us5pMApy8egfb6cLw4l5W8tBQ5K1S+40yFT6c
bl5tTQWpZVUeYuAMMknIbKII3G/xpEqu2LqWSNu401ErJtHI2hSBoC0CNro8C6DyZ5I0sr4BiK86
7YvhjvJkauuqgPURnZdlWZmwnQsJKxEDx9ysXGNUTdW9q0Af+PfqKq0ooW9tS2jKKy28RQJOHNjq
jqcO6xUKAdFmmwBU8ntoJDtL5O5SE4VOwiFJ9s82swYIS1B/nSADRz1IvNNZcreQSArkoKyc4Ba8
64/31asgkGOJSAjhekAxhThOk+RozN0j+dZArcEQ/7GJf2Bos+uj99dQp1p/1twP/h7buMyTkVse
oMdbYUXhmw20KScfj43qcZLZDpvsktOHHhJgHoxXnHgGxte44Gbc4d4stUEvh+ZzNYjSefUzHMUW
Q7wrXjL0qEH3exX85W1QRuY3ReUoWnLHQhkL8tgrqYoaKrBtEUvkV/JU3OB6GnzeiK626ZJzijhx
cO8vLltZhCQ1+RFhJoLx95VUpAUt4TPl4xFSKAtphHwof0vr02+KIRCUT/ZGp54QWF+5eRd9VZGX
mUb3gdT2t7CxDH4WiCs4lKm/aYDqPh1dZDuiBsxYo3nb4dxCvwUw7iI9WwDLlLA6FxbO4oLqmfVJ
oOGMrudlVkl52rV6h4oFzejSLui2LFmi2CjEImhdHzTMH2hsYZG320yQfV0X1X2fxghx5HDMclAi
bsrhH/QYMiOLzXvI+QF7dj608YxLduv+Y4hFMcbdem4RVuq4KaxwXFrFLxmAptK8kv0idJntJr9x
Kn3XBgdp2HSQhAAi8S8c2YVGXuG8ZNP7y0du1jkEh+Tf3/rZAap8mpth9NJggvQn/WBMJopNSkgG
N074zW/UQ9MhQ3DvJjX4V8adzeyaluEUdADbFcuZC9fR4mufY2SFXR7yZW7t6EfmIlFkWMOJ+gZq
hAhkVWxq0IQ1N/FisQ/tyQGRPpWnoTSBmdoaer4JWruZbvDB3jZw+9uPUQlFTZZBBJcwcHgA9SyJ
L+Tf7lmjNJtED1l9iXHe0ZogDk4Y8JtqhuFDo5dcTWzH+AxMA8iInMMU4B8uPi8oFBAu6xBdStjI
JL9ZHoHP9ZYtyfqYwa/5iKCaS8thRyqjN9Da7UVv9Zu3NAnYb5okuaL2FL1ec/Yhsz4g9b03AwOk
5Ho2Qvtn/sJLjpdCHXi8S+fgO4ZujrLMrG46UJPZDjMPagbr8YbV+Ne+C0UjMLiMy4vSKqB4jJKv
ZBMWWiUdiUmaAa0pWTARhf41LzkV4UeOOPx37iLAy5GrU1XO3stR/5XHReRNpaOQHLQFL75eyWcG
dXUPyAtLJKw+ITVkzxgKD+2W8WIs8XqJWBPCgu96Oo9yibg2CwJCU0hWjSTMyEJUdPhInO0okXtE
Fmj8yP3kBPTonQpGI0OiQ6SXK9nul0TX4mDJMxlm+iGYtjNlXJdnuffjeoBRIT7rKRUx0qzPpBkx
oZ3TEvSt8k5qu0J8m5wM+ur0aHW2vM4psZzwKwSlKtNXRyT80ay94MkFxoMPN0eg19oF+C4MWgfm
s6RMOad9BvQCz90zRPUOWnZUUF76ESU+e3G2E0cOO4oy7c7TNa2C01I2FX0K89VvOtjjXJY23Cel
F5bLsz5iFxXRW92PhRKKiN0fAt7YY0cElyqUyQD3JDahXsSY9hUtGZsWcsieqJW+iOY1frtByKRu
DQulpteDtcT1wDjWgWECW+VsAiE/Q7tJ++vgYTpgN8JC7CuYc3w9P31ktY+A72AJ6PuaibL0YPRF
MdtiKpt5lNv22/IFwL+HCkXwJKqN6nTv1DFauDEjf+DqfLhummt7VUU8gdLh03WUa1FIqtQEAvPq
mB2IuCN1LsctLAMLByMtZoO75wMG9o/B62/yEca7QhRVhV+lASv/6qT5Opn7Xib1BR918lYamYRb
qFX2QnEyca3pqgo2w82Z3wH0nGYhftQN0eVRpkzI/hTKkqppzn8Hm/W1WIYpJTtDe6QQ8mo/LUeU
IYDxke3l8ul+dS5vfYv4alHDXW0UqILeQmccYd2lc2tPuEgyPLbKUg015t2Ww/z4hsYtdzj5PyEb
L8VJmobgm9gGFy+wZ+tykR3Kh4ZoJBysZ7wmxEnXxHYwfSJCl9054MjnB8T5hp1JSi3HbOW3V+lT
FiZ7MLbFsfHALXttWWAsOFwKLcqqZCKf02qAVUq+UBpkaVSAaPBveAdhYbVivBT9jjHIkENIZesj
NVMtjmkvCvs8Lg2+PY2DUNn7C3Oe0szd1Ol4KvxePylgBmvgfBkskGWY452T00piYZaC08E7WXUx
FfFsnvQDLGMJYmaMxYbHJvH7pEnuMKv8YdqIaul5v4/AChFMiC26tajhQRICXd6H7sUzXaYNjjEe
/HYnkqvzw+RnOeHzu1n7VpRP6qh/HdwOtDWPccev97KGvUSSA5FguOBoe2QUSV/Bbi0dsPoNptZW
2YOkOenSKYk71bcUFm+MKXNL16+FKsjc8sFUvqJy1l0TNVS5tshI7QRoratnKgh08kSkVsQgvD8q
SIW8uOGR/9AJHxl+GifSlHEVwmz0UlMsg6lxpTGz0EM2ybcg6O1kFeRvsb+pPwbik+mShy9OKAuA
LN1Fu+4lt7ZOUknpWvuLQXAHkul1FA57bpB3Vc7qTWsBk9haDoy6MIsBwuY0+IftwhG6rKTabCvB
thR6AGP9K4kIDX9NShNn0zF3o4w842S2VvY2D1ZI5AP74NPfksPPr/lyOwJaDOPjMKoZSW7CwQrk
x2BLZ1PoW3J5JPjEyRoGJ+GwtfHIu6t3Bb1xHMwU8vWhTtKgtyNdyHNWMKGwtajBTcH/r0CRO283
CYi8X0i1WaCJFHgeBC5aHY9JB5zHbNLgTzZAob9pnKNmMD9H0HrHNar07QDPxqyhD+IeNGA9QKCQ
HngpGLIRlMo0ewzuqA7p7MKjssSHTaImVaSaIjAMCZtOQeFTTNoY1+wf2t5OKRRrkqhcTbPaQVst
K/abp0vXZx1JKs70UL5N1TQJhGzRHdAn9eZpTPg18XG+b2/TJq5Ki8YQn6CKjD8cVBLh+mkWZdVu
AZDNtqpBZr4CXiL384/LxsBNs57i7iGqQNtsti92gd1HJfvh0/NuEr2mRxIAnkmszYE5QxRJPW6e
D4azevFP/FE5CBKMw/649OcwXb7YmdWd5geaEI/w5+S4oOHYvIC3v1d9f+C/5LJW1m2tWIpexhUS
g4LjqwLbl5H21eXaRxcbZFbdha+LU9OFaaWk5fXOP9zW+HOyrAdM4MYABHAL+JQeLqKNT/UK5FMS
XHQAg0Vtf0kHySwSZDYzAkxz4JJAOqp4QNY+3iRElBQWF+PEGl+iVk965oFSZKDblc0NXHokM6/J
pBsdFA1MMh/Pucmm/KdCUwdNxdffIuwutLsMKLKu3xcJDfdTWrL8ikLCIrYDsgDC34eBGxapIRK6
c/CltJXPXpdryhr7o8Vp/eMphISQPQwSUq/kSt4mNE/xEENlegI468EZbHnpBNpw73ZOwrlwjMr+
YcpMZYTb6pt6elK6AGPJNSjsBQ8dHRxg1GBr4iZFfLUsfS0ljGVLXLSiAGIAMlpGMI1ZMBedexIe
2i/HEGOifHA3xAq2hKTRW9aInxdJdRZe7rviV33HgkAmUdNzVgyCCKw2knAJjybu/zI+4gB3nyzY
IYZR8JnWlpn20ipoiJG/p+QMD2udptedK649babovysHf1nocZjSvDtj88BKfBqCa4Kstx6axMYC
WG/kjEhH7ngJNtPkCLe3NBIVoNoQkQXi3Vn7sH0InxRBhJsIx4TOFzRpf5hNbfzDQfkhTHxvj3e8
FbuGHyk1JyldFlCrD/VIVejDrw6k+hvxuqlLU+Ys+adgHi55jAPEGmHDqdNRLf8abbWCEUqARTB9
pfbPnJvvS4XGYneWpSaoqQmWplalLl+mLOubDZ814Jq5U3GpA5ld7gRNwzJGRb9YZAILBjRucrlV
MXOJm0lx233AVk5M/he87QXdFvrPVN1dpH3zBhn4YXf5bs9BCOrCiNYH5YcjhxDL4cxEOWGeS4f/
niNUDNmWeA65TRccZAVHBCMMWFjVHu17E6D1dICmDH+RehS908W7XxDvy6zUt0xhFxv7E2Ecbmxk
ejekkYMQkn5UBGJuRucekWOTsA5r71EjxiAM/wtgEYK2twlKzxqpjpl6V4y4EmPaz7RAwI3kMAAw
9XWt9tZOZzQgqufOhizQkJvIMJEWJs0idZCcLaiU6/XW+dzFuNUYbagS8bIguvfLdTJYP08fDXrT
tqtf4aXWTFoUweLl/J3qnHkXHIZPhpZZkRxcuGeWJdEbwUcHro8HZIzOLed4tiNTe5TGvkOTVzE3
3HBpdQbQpGgho9oSEvGk1DHziuxxr+5kC7UaGglteUQ24IuwXHtrz3FydYgNpWu4/NCCKMHelc0a
RR1wGiRo7xNpdW0xbG8AORwm16WVdPYwkWB1OPgLM91D1Q4U8AcHA5OjBopXtwBFIiIesqNH7SBX
NwEflM8ARDe8IQ8tOiLvloEy+nVCjv4ymUccRHKg9CPLa9s2gVcWNVHlMPmD0cMC7F8yMAwKCfdu
3yjc30bxX3sDN5mIIoGdADXA66i+VFp/8yLKRK1wOJizh7axnFjhB1y5jlTRWMCEmOg6oZbROBUz
8ClmjkzOsh0P8QZHFHM2sA6gwQ2HBtb13qCF8wBhFMm7+YWHL/MemZ86zc4DE86JC47fkpSPpDd+
MCi4u+1ISL2vGlJ27onADdBB1bvciCISVzmyRbGlLX2U4Oe9z24rOQFtGc7idAxY/6a8JyPH5udK
U/x3oKC5ZkYmb8u4XA0RZVtvATjf6H5oZD8kZs8z42Vs3buC7Kn9GWkrSIArsu0XKOKmo2JBKsaG
BMzxkSOYNoqC9TU4TGngmLQobzPj4ppgQl45IBihB6Bt70ENYyANskvkGlaJdBGMoqsBgVn/V3ds
qz5ivLcNrcQcgEgeo7C/R1mc+khOo4/QcsyzQ4nI3TKYlcmmpEorm6OzqLDN61BqpdVZuway51HQ
63rGYDjD+37RMjsbGBBdltnPR0hPgvE9ngVixKfQ4mSYsJwkcDjOtogUvY6lER3NNXZgkhlGhEzN
JQsIIm7tCWA4yIIHIoWHpwBooDb47kmgTtTZW4SkO/PWS0l7AH4Q/8P6+P211e2Cz7FV7pd1LF+M
xJGo3Mxet55zx7yXbWYHOsWZski+g/4xsmSBZLGICgeqDmPzxKZjiSiiyysUoAUuog3GT6Qjcruh
6OR5troOCvbDn69Z8pY86k84qaZlhloHIdW/Iv6LciDuQNfb00KlSAecqeC6iuedyxGpatwOVgKm
xxlRly4rIuKcOYR8Yks5Hic0hBsruc8VWKECijrll9Fse8X8TiErBQVjiCw3bkZXKL/FtFKJr7AK
igNLmIRjl+MZ7hVGduXBvbh/B9URyqpD4NosltoqrAEbXd4E3+hvuGZsdlbx1Es4yBEIS8oSUmMJ
pvJrPQvSWwmMqBTNurEz0lqdDfwE/PXoB5n1+A2ZEpbtjkumGX5NP0GHdktbtFCRHEaJzDpyeb8G
aD0XQoV2F6V5PywbEMdBc/6f8ZN3VWRsUKb96RhHDpzCcJSYoggkR1BjJTnq/SAxwjkPRJV+FFlV
X7w+F2/9P2jxGSbX6yXnpSuHofp63/K39GBKRrqz9TJZyTmjK53pQ7AMMkkfme6R0hImY4tWQYHk
xmgDbQPbEQfK3YtTZngmCbDGaXk8qWM8tR5qzDDuztCK1WiH/hTjEmkMp9oBdTdsWEqABvn8+hXu
Mibyx29tvsntcQX80zRb1NW1wRe8RMqw4fVtjobzurFEWtWdbdw1oXv9dRqoeKEsTQ1UfMc0R4wu
70gPWtJ4oOTQqE2UmauiN59m9qbBSO9QxEflyTKFrGF3o+U1R/HP+it1RAAKgxl2rc3nWP9UnJI8
nOBtBpFTNeQoCxZgMIalEGLD4FgvpjuubbWq71XyPMTJ+QdJgglBJw1HDZRklnVJRDYGv0JjaweP
6+fUFR76PXfbLf0htPa/cp1D9V52hEZEz9wsPSF4xe0mFcd7Uur+W9KjdogHmkrFcSs9tK3df6JP
8M5mmF3Gm7REf/RxNQFRgd5i9NmU5UliQjom/1wyBgywPCE74YzXbdJHQYWOwf9YXlrttsyWpeEH
vqpIckDky/c7HkuT1BN+GblSfCDXmpStQtqRT8MY5CAU5nOHRleK+Xtr+CG5u4M+FSmaZ5vA7qw8
DiirEgMAGvSFKA25TiS/Z0g2if/ByNYlOmvfaL3x/5zxt4nym8tMqSqIA7BS6Uw3Nl8CGg7zuEZ6
bcMBFpl+8g9ftDHBUg+wAb9CK4JGY9dJTixmK/WG98P5FL5MYM4ZY5HfLc2PPtz0XE9EQm6bbHiL
9ujEt04bAIlVRsUUWzAT7DLYlLXGkx0Vhy3SMHWYE8GTVUPUmxleY9KDwCZET+AK1awnbgQ/IPAd
UqhhmFt7q6tSYnL7N6wojkRX+OEj6A2VbzxvAKWasFtSshCsS27cMo0IXi5qalw/Wed1xNf5LXL4
CCgZrHuf2sGG7SnJPIyPoCmIBRmLABG3nrLgIhGyGiDSV7VO5sqpAaqmgfXN2W5QXHr5caSaO0JQ
/J9wOgQqH5JNCcODl6Yr30FFhbtt1Et3dzwKk05kQQe1SfmJGmHzc48+V/XQqn9teYS34CQ0AcND
d1hDWMkySYqGvZzC52K/zw4hWOlYy81KRQ8rLjfWQrXqps0yRzkQ5fxc63G+1SOBrLgQ0xuo+Ruw
S5PwP7oKQ5sugdsYH3h47wxVGQdQErjlM8lmVZbPKAs/6SgWE8KxAETmbMAPb7YBTfEiIE5Z/dtq
6ZK6PdRo23PY4MlD92PRYcJPKgMJYywG5XfUKiiKlb6gq5XMS5uibeLvob0eqGSyR5Gd4behzlqx
2GdjTd5pxubflOR19DcIwZ51LqfwW7oPCMwjVSETPMfm66lRth4mt0n6EgDlTJmC/pWsumpoLEl/
eJwsa0ExfMX+AXFnUoNfLCeVktr2y1+/6TDIJO9UMp7GXGQNQ6QJnGNUBxAJKjptEVY0Qs8LXgZ1
/BVYtyRh/p9DRvOaYDjYQd2uLcb/bLH2y06A0VJhqKTySsHXhWzXrEu9BU2oMqSNqYHFd8WRQQSl
eVrHop19+SE75J411NP8dgCnz/QTLfEbFyOKZUZPhHtb30mZ8rWz5r5iqkjTwiDDmA6hAimTebyh
63ir9blI3iVfZhAIT5mhK1DUN2pFufSTPkg+i/uwehkGgN+a+vFiizNyJhtlEIwbPE070m1rfHOi
FlXMq8E1apSAqKgR7YsukBCjUnmbMIHx6Q1oGL7jtmFvnV+cr/AE9OvjkLL8bBuE0aWdTBpUE8NL
BQMis/l+TpDPQJpxO6NXFZPSPgO3apKNIC7CBM9V9561UX7DelZJdDMbtVeUyWqTzRmiUHtjd78m
xrbredz/gZx9go08BCq2pdym6nchf7VMRxWnWDoMYj9VWHqwwlt3jnhitky1dGTF/q9rWFEAg5rl
mi5zHzCqwpgY3nNczIhTpjOIwYmJtfguCffsfXPS0tbIhHyTrTDRLVqf61Isuvq0kFXdpdzJ8N3N
qQxmjiSVwzslfVWFUQ8/IENNzOMybJrFiMCU0+gJN+B/un9sgjeWaBSutT+MrQDSnoCnj1jJ3gBO
uIZSuvIzmfxd2+d4//O2k+ycmX+PZS/1XMvmAo6IIJiMZKOW2qsM2hJ2yi8w7YetvSTMtdk9BCNG
uoqbWhno+KmvDPnh2eN5dfhs4ChMKXAhbEB+qLoSF6bbaXlxqCRdbAstLWnDoSDjjv3VAknNtROz
rJSrFGE5ihpPyIkXUcFKRSVbEA7+HzdZN1AU44OAL+++RKnoatJts5OoCxFFo/5V4XxjFbisDHHk
IwVI4mpZwzKmzwou/Jxl3DAb0NI4BCEKGWjlVp1AMfO9ueJiHjPnFD6hVJ/yGQxVbYJPSWn6Cilw
Lc7MByHapJi/eKaij17j7ltLQ/Khq4xFiSQF/2v4HufZJn65Yx3Rh/bm8JX2l94bhqToBqRLiM6q
r70w4qKZIrd0EJxH5bLYhCVBRUR2Q5pNzrv6JPNevamUV2p4SJLNBIGOd3BSrjDOMCvYOXUEluaD
c4Toxq19LhXphCxGAcvQ++RcuHu3xkKGYYD7+12RLPpJ4Spxi1ONTYOsKSUuB74CIUd7gPwpAPd+
HdEg13ZRP/Adx/ZEYe8D/8S8i8mXewuDu+skWhwm6XRzo/nt0eAfWuszPk7c135XQSx+rBDDdOEC
cBGTFby9prcnB2fsVZQ203Z+UdtYGj0U9kmt5T/1Jw3U1tUne1TdgjcJrtn2qGMaM/eAKxKoJtoF
cFa/w8ddozG/3JzrV2u4OjF+VGvelCJsl22Z9vynNi3y1k0hPKrrQhA93GAiJynm8Ma1vhRBwcfo
V1Y4oYVk8f0mVIV5j0uNQsJYD7PAGNpU4rrxhHLc1jy2tATGPGWVTC83/Dmn84cK7x8bghtjcyrT
ZoDAon8GJKlGHoOZBJdUrJ23VMDi+13Hez6hmfMA/0Tz/bDZu2H3S7TfncUS3+iWaaYxJ+AGrkUP
+9Qx2oYOR5g0tPsxOGm/DQXBm9mVFjEjLEbdYh5OHC6urikJifWEhdO7TO+wJlXPuN0suN1S1StK
Fr9hRjcsCzj9+PNwcBkHlfZbBLbWNe2Fl0oPJuauGx11jbblfdd4RadupehqPoIqm0COTeb+S22t
5P7L2jhqiVbv2fdL5+u0jroo8rNjjLRydAdrj5kMa/MVdw68KVWoguCz+1N+5yDyOYe0jMSVlzZJ
dPhXT9CwJg3P0I9wsu4AS81I2dBEalV5t2NfA2xkiFP5HwXfTxkn3GKEgWF1RKffNfO3uKlakeFB
MdhuixDp5KWPFAjEW0h7IQKGmQ1UEuRwiy2dLKgYmtJeS7Ckr6rm+uCeZndwu9Ed+qHi3jjIqw8j
LKPrYAYx/wv+prfI8St45famQWKQUhjjXds5P2TBM40ky7MQf/4BK2JFKdb4RkwCWI0xTBIzZB/6
IQ17pP2YjjGBHCym4+/vsdMkQajXWpMtqnHR5HzkEShVDvEHaA45fNNR+Jmo7Pexl8t0Itzt4XOu
oY1CP02GMIxs8scS8HDiot1int2pobe6WNtrOvOVK+XE7/m6Aw56Bc3E0XnJR3J3lIQBLVoeK7VE
DH1hH7x/b0aZMj9tsfijWyaHw3h70pie1MedwVpIacCXkUEfJzO85rXDFwJy++SQfacx/+4+Brc+
uw8oEX2gDQgSikjWZYxHHm3oOX5FhwTtzqQystFgFRPjfeZGHV2hIBqsWr52UHx0RGaqXue+DzP4
sL5YztYKtnUxj+ArC3N4YQbIQxCC2LTfvjDoqDb3SowY6VwJUHQmiFYRgNkaof1B674fGMbjosgl
JTCpzDdSII1NqeHG4IA35G+UQ4rvJ3235Yq2JjC50D8j3eR7zJy2+qYfUioiSahuq7/uUAXoFgcb
Gvn5WVvVJAh4mhFRNiyGnqNUzGKE+vbX/Su3g/CJyhvWmiNyDRPJ5zbwAQ4e2tESxG+CAc5qD+Z3
TcB6gZSUpuC127oRTEacVboTZCVHM+e6GZmeIqN/mekfPo8W9QuYbMxQjJ5593nhjaX66RHAREhi
Me1fvM6/6iZIb95dF44+SvejHXrngU/aQN6moEoc8wGYuePA9G+cMp+AGldS9ZQx4vmSimKtB3io
CP0vVHxUnQ8X9KQfI6Zmk9ewSDsc52xfLVDC8Top0zMupS5LR1jeEiMVxChNxz1rX7AHBxxstE0o
/G/IvgWqsYza9JajGugBdeI+qGpe2HdGTvpsxluUGRs6pMmwPga/yYL3doHNkUNwli2jNAkd3c0l
XI7AYuKzWowOqKEcz+8MaltRvw0YgSUUvBuAuUaXfnj8mlT68JpE22KElsbfcmnVALt8ZN1w6k1J
MSSLtZjkIG9q+3UXc0dI5PckaIrLGDYR2K/0RnqQtqCP+eCc6D7xSGNuPqaUiqYb1VqxfSRY9Yl7
/IJymHGtB1/seDPuuP3r1LkHNXWzwQTP7bDpPa1d315wEvRLosA/H2lqapOGjaDmdfV7rQNG6ATz
yH2i2d/6e6rbjd9Rn0HQSObx2wNBp7pxd/wyImyIUp2TYDzH/tK988Ygp/mZsWT160ZcTuocT3w0
j9R1XbvsARxkk5GzKsUIocsoLl+b8exxeYRZHZz9VQBjY43AEvRG2/EIkvPswrmWrs+lucT2LCzw
LhNDhfQOugDQ7pLhNEo5wMiOAyW0KMTPr7XZdNwu949V+0bXHadnKPzpJANleqcGW9DfYeJ1hsW+
ei/6YA+SKSShnc2e9WssMaohmUkCH29x5UT7qIE2TURJgnydo314/CR4i6+YAn5zAmVJbb07LdM6
Pw2ZNBOsKbRxMNcv2pfFmkoPqwksCzvLEi3isFjwgB+DQlUpR/9swkmyXU5vP4nhTScfjQeGeYt7
Lp9UBxKwYy1NTDFGh8o7QOXC4nRJy1r3Y/UDXhKl3oUGi/2tAu8gxsgVCjEjuaDRwr3eRQoi7gQD
1pK4RZm84hA8AQ//DJigbFGMzpFzsdV/GjnAUd0xjnflj0/7/mMg5wYdIJ/u81M3M+j5dZvQZ8xL
Q2aVHmrm1CXuG+ycWQ/MeX9s78M5eMcFpuNqZ2YepR36Z7b3d9M7q0xJ/3TiXhbN7A20N4CqDqgl
8NpV899NsKZbmYlmYIC9JriIGfu+7F2P3LFLB03mVNumJ1omDWvExyAGLhWhjHx9XEXyv9K2pXeI
pBmEv84neddG8k/M+U6xCFso6sv+L/Q3jJB48gPixtKEBqo9VIXU0/Q1zzy/goOROtVdzhhpZFHm
Ilye6KY/ZF5TsAHS42tb29atrwcg4yx0lP5J3LSQjEvIwi4jjQ9k11rR56QOEEuYoJ1TkPZz4byd
F+e8ppxrzcjz9VMDB/pTSMOQvp3ZtagbhB7ai5E7k/vORW5tf5tgudiB9U8Cg8CO7+friRHABYds
+3K1nlFhKGskBaPBNU+71hcQPfH2Jsgk3CMc0llnbVZdLORdcTVu0qNIapcsevmZZnDD6P0wZ5Tm
EOK4nA5fcOm7HoI1futwFJVTmB/8kbajOpyq6UKHZfFD5FIadcykrSpHcbpiEKE6kYG5bi+mr9SH
YU1Ybd01czJi+L6tkRecr5Gg7tBvLneBxqsS86n6Kh3Em3HK/gXKm1bzUT84zdQpv6cLu2LEdNKb
6DrAnUljCWbp8NO5aZsQtUXNmwfdMjjhckLVySMF3mwOPUDuco2uS4f9ldqj0ZZSL30n4zSQkSJS
ZK0Nh4ohGzUP7IjJlQKVYg3DYttsp4OS1iztTSbTRvH6FlwuqS6lajCAPhY8rW++nPKZg6AHm+03
YuDdafvPNMB2Ei59V0zDV13DHBj1HXO06+YLF/kgjul2FDMFlzI4OhtXDcpsrLadCz4FtOX2O6v8
EpOT+6dNtrFaa+tdq7Wv8aFvTD+bCH2s9COOQiVk3j+JPm3RUwaaeFbbHzjE0hbwvVPtHkHmDHXi
D+iyPicq46UE40qojIvzvDDN/RsuAilKR+d7U52xmDDVZVjv/qBStL0vkcso+Z3DklhqAdQ0/8R0
Acn4/gafV7o5QWqBClHQKmDtYYWM6v2XaAJpf1Gyb+WbmgA/vvx49n3F9R7VZcSuxfLJ32R84r7J
Iko+Tn44rYMv63Xfg2YKkpjO14Q3sXUHvXhmaCbLQ4Uu71oYeTgAUTwCRDSWx1TaP3Cv6hjVNyHc
9/50p8HqZRZh5N5gUgQ9Rn2s8X2BsNTbhAUjTmFq4J1C9lfTjHPvT5qRcWopP17/5Ywd/o8+WRWn
drb+0gkRX4BdaYUuTtFGfCyy8Z0cI3pQuP/EgfLJaLuE4FQWQxTcIoj3bsnhR2oAMxHNjHdNK7HE
hdXzrNFp1saVjxC+w5GBZlYylQxPbb88SllJqakrNH7gyWdpeICCzFwN06E1bYNrwj6mIW8IgMfC
VZjZOuDEpxshLJLxZ2zavumqA6xT5sJCaWGszusy1GMe4KakhDnfuCSbY+VeFcCQP9PqdCY3P23U
44V7oJLPa8y+7O5SCSvTFr8BCjaxwFXtbWAFXY7MQZ96kzqnaZAxECbs9iQ/e/HkvMKztzcRlzo0
aOG9tPGHfvcBF3UKwCfa7s1dzGEM6tbI9z8Z2w6sdNvARFClJM0KiZG1vmJ7407+HyMCVva94zdT
s7mkGb6K2bcQLBVpwE6f/foRFEGfpswSV5qDRllCZgYundqxy335jZT4uuGVtfTJvOB/RczHXwtn
vMFXplQYJ6FHGx5Tyh36ThFxVioAHqKu7q6wVFbvtHWQDlXUdDyl3LY6P+p4GWDUq/ZwZ0Mi7CzO
t4JM6g5vYb5FpsU4SOqrse7/MisPTsWjI5lPVXI3o4/3PI+4afQQ8f7XdYzbgttUlv9pf6pbUBqX
6eWkPoMfj5ECJZwvlrQnTku5uWPQNr8DwZbRLJi2eZ2hcCMgN3B89XF+/mHrgtuwVZLmT+7OKGDH
r75SP8ibVB9UeYMNVgzSv6dzk1xwkUBtfMniMd+u9vjzKHvaNuls+UdxP6jUBmPwpb58NECwlU9y
s45bf7iiG3G/scRQZflQmZ0+43l4sa0RPV3KQFa6tmhZ4ifDVsIn9VNSH2ev0A7svSgXHuOT5eKn
Otg6mIaWj0y6PiWE3aaTiMd8JyybMciJx5WnGlwBcVx/XPnvE6+MzHnLcJnwat1blrvuzmobzJKl
B8P7qImjksA0LFZVuEgbWTGe0WHcd0A1b6Dh7W6S7Ij54C0lMeLJ8BNSG84yGZmEUL07yyOS2mEE
qvZcJdqEXqilbsaPOrsETSm0WY36HNBYucyYuUoBSU5mUujbWiccQ3zWAO5RVwz+B9W25jAVm35w
pMO9h1YqOZwdGF3Yd1KCEBkhqOj4Uqo9XGoc1ZWZeWGklw6XlIes8ebbJzUHX9xSjRQ+jMkD7sKz
B3bvTAolYslCVTx7wQ+rr5cO+9MyEgKJ7RpZGm/BmN8YIuqlLjGiSxL8IZGZ5oWsP9d5yuKuK1a5
jtd2W+5q2vQE/koYPwecoM3LzpxLfJiP9s52fupBhFs4KPMqKc85XRSk46a/JCjXgpjHCtrvWg69
bJHAekq+Go+VtsY8F6BcSzs82krXW5APL1AEq14c0ytJ0Xk00mKj+whGVRXdT74/5kic2bOWfI8k
/wHbPvwXfFwFjrxn58ShsF9f3GCOKCMu7M6zPFeN0MSx1RXRDX7ECm4JC78LYZsuVO9cXeV5LG9r
xs89XnHIlV0fXnAnoLLR9jM/F5NT2VG6paSWcwY1RPcHG/R6QDdDS5rcnWjxHLqzbtkXvmZLChd2
2AUHTpJXceRv0FeFJlcwebHul7TNnrdKFQiqyFOnrApw4VKFro9qRPRHlZn0gbQu7j4qCkIMm342
sJ6OLFDr6u7V5DdNaoqoZnTzwtpQFOujsudSjhsrUPGyVqPH6rvqkLlR4QJwIRrah8q6Fi7Ec7nS
MKIVVxgM0DR7oN8M4QvLjQXDGP3lyhWoelegu7plH2CQdVvsPWg7qBAzPFIiA3eXo+nNFIRlxnpS
J5hjXINg8umB/dBuxlnxlZIw+MU5Es2nRTq7Le2KzRuntEvi2YI32CDTm6nkEbJHBpQTkj0x9zFw
Kn6UOrfNSZD7I6rrPQu4vLEpgJ1zs/VtFvxCp/utr80uIwXlLurJ8DLpZ1sQRJO5NJd4QFW9kHMi
94diXtvwC0UB6YzzAOQmS6GByFoL3Ga3v3DCAKadgpiUKfOXKj/ay/AgUfxzd34K0YB9KdtYjD5u
mKtn+AASP1hQKYgLXGqg+iv0BauIuoPEF3t/nroM8+/8NDKOpezC6RW7iY2OeIFCiZSP5NfXyiBx
nEwLpXYn/0qA0oJLxaXu08eZhInrL1w04uxRPYSg59/6yDgkAA/AhzNGMygQIPntbT9M2d4dGVRJ
2UERINX9SSHKrnW5aAPdp0UjweQY+yfKhSbxiIKIuJx9hT49QlYtLnJMuttN0qCfppkJs2jl1oPb
LD+ZEGuwxqL8v4yVn0Yob6ASwYVQBg8AKtyIc3z9mif1sWSnu16UhaYji5mJvpcwiLFjFQ/Sp/0I
8+NjsXDELQCBDqotIVCHv/Es8i38Vrj/RGyeW6IAn9tvw9MWv778fEcOA9U63gdfURGKTYHgQozJ
jJupTtrkeB+Ohwh7a+jt+Z//Ay3eZX1lX6CtYVzTXCsrwC6jhly6LK3pQKTrWOY+Z9MzGRodqsdM
+i5zlyZm2v6c3ZPyGJgwly49PhUJ6ND57O4IwaMGPWhsF4RLCYkL46darF1dtfknQqxuv/0bnL6A
uKKbrFYW1lArBOYhoUaEDAVv4+JNrVmVblQ/50GPPP0wz4MafEW7Zsx/CApiMAAjzjzFFNLYk27g
a2LodwTlKJ1v2GAL/J3hb2RNOWi82lB6qj7zzwvfp2CpZGGg/SOK/qfq6NT6N+ku/R54E3bYwm/H
HGJ1DOWDqcSk/IZqF2BkkdTfgAafCUTLWJei0HLeRBHd8T3AMzv8OLAIieO3MpDBDqaRcBZ/d4OC
ULCBH4yDs4zcAvKwKEY0LAP/bjngfdOMKPgT/iTz355MNR1T1sGaJU233MHPbhR26URbggttFdFI
e+qb5ZD4INr6ycDMaQZ9oDCeQeNSl7ZklMkv5D1BLBT17Pb+Er73BNUIkHGbnjvDwHp21sZSc9PI
/qzdggYArfqhJX5v8dXbquVvV3dC4PtGVetkr8HRMt8hmSrV7DzdtZmTL4R/7bCGnsEJw91DXr8t
uWVT7mhEMl6Oa/7WK9Aj51GhTkMKrO2srSe7yYI8081U5L5pYumlLpoMy1mDgF7omr7Ch4+gRSVn
aFlNlNcIqksj+X9g1LLDOROmexx5BYix8xFcrhFgmLO+VTwaXCBVrgFSpcDGdzWreKD9sFsIRpsy
+Gyql/jXwErxlp98hL4iqi+tl4LMYiOjpDNrvRgKPoIMCg6pTbH/yXfYcd0albv2vp9s0dmwuv06
FsCJCGVtbUr6hotusVlnthWB4XIL6Q9eHDkc7FJ+1ErBPCeEECLCxtI38urjNq+SsR/HBpkZooEI
hLpjuAbJ+uGLENZqCarT6A9CAHw9C3n/sQmI9kHGdBZ0LJkSLW/lep18WoLYPzEwE2I/to4oxOTO
b95Mui3oj8RoWKvKehB9pkE0sFiV+SDWXBvGbvGS6gf27mz1+fUYLHJldmAhB/paHW4itOT1XQQ4
8D9z+dWvzGPsVKkd0B7J5Y+hUgluFr9yH5x6GdmgCjDZ79QIh7pa3WvpNPm1AUvAocPI0H4mStOt
HpTCqxPhsd1JGQhVLEBLFKkp3tJ9CICf5S2+1l2Y27uo/DNSdehlRF5sKWWFl7kbh/rTqmIJpSG6
ku6G784YU9r+jdvt5MTlQXuYQzr3vyeMLQyBJcEk09Hv1xt0254vhluXci8YIBt8G//MGDB6ol0X
ghUyJDdMHFowItsSDBQtrz7lw/VRXSAkOOOD/saKmpQ4v1GwHq4y6syzBpU5/tEJu8w2Bsc+h+LC
20g1YBF1xCLQQ13eaHLqhkKW6uztZRdmyfRNeAAmwZYWxTnQRenl3zwT0umtOd/BNgSSmpDBvrO/
qKmMb2ofSc1692QeL0aBWNDxNVA5jVz5ywIJwzmyub9UelXCC1wdndqrefV9tvWmGfcjMOnX6xWs
b33wEF/PL2ak9GhX0b5IjkTLRpT0L5EXhJ6gufEa1tjhSCIAAiW3RM48SQDurchJAuQwlaKW4Y5A
T394cjO0T+U38KoKENTQYLBSeLrvdyyFhD1NacKh5t5b7UOLwop8V/GdfoiMAfQ0NkpwFru+MdHa
e69Riu4tSPU92KjDwcDu7wh4HqpJ3ZjpjHzP4Lvb11+tBUcjRxhJHj4pfK0QLtpgWB8SAOgYu3ha
Zl8dzn9oN192FzAlJy5dhZu3oi+JmTJe3n/UT4fkET2qKZjwfX2N+LO86XdGoavkXMRI/fYM/wqO
ZBMHHyqKqZR0JHkid0SnKgb4lFDcJlsBKuJyurJ/dab+AhdApzE8jqhdKsGZSyMQh6xTYZQEZ0yb
bkniEhdBeufWKaUHRcb2JZBuqqFzPHadVhTfDohmVuC6RvOukTK3SrE75xDWULbJhNWMoFkzcw0x
SbsSqsWWGtMTmR9ZC9YGRAzSbGYgh+dRDIrXwgI8gwsMjw6gJBR0ypSgMugCrzaQCUAnkyDnlTFH
gILSPYm2xxmMV/I1+RW5QVO3+ZgzLe4/Eiq0PkAr0voOOmVrzPk+R+r3bPp/aPP2iHyq7zRc2apn
SV2/HPW/PRcCHk6xV6hIQek+9Ua9JjuJgXW3dJo83Ro86UHQL0koshYqS2sXCI9g5udhNvoCjNA2
pmM+m/TBparuBgbuicCm3KYLkj6yojuKr1WQxwF8EEz0bBJFUPmFpRsgidouuQYGWaD2Cqa6y1LW
mKfU7ZQtOxzuH3s26qtBCOf6vvqV0ocBwDIRld5K7KnbMB8f8Yh586t68mRWaBrxdUnc5BZ07HXM
Ufc1kkDyOx9VI43WsBs47zttx2ncgqWASw+mJEwZ+kc1LGqrQBo8G3WCGS8/3mvLq30UxKi3y/Gy
Er7lQXfxmakIP7IQXE0RwTLIX/HkHBOf3gR5RQDjoC8eQLWJN7wssB5wOjVfwL2F2Mfcptl4hkFg
fIK00MJ+/q3lgkNP5nWOJ+0lZlCT/kVThG8SSi5wOAszSYD7PgcNiOXsFBA+4F1SYKhqnUeW0jMr
G20cKXDFGgzKWtapzbx0/KiZn69QmAKyY9jk6uHA4svdRc9H9bMBlPh2TJ5wXsnvykdnyVKtDYB3
S1txheqA7p9dPVIvi7T//IF8y5l1+wiGnAwF9045dyiBL8uN5TJUYjEbp385FLrDZHnRIotaP4O1
SA4WbzgSW6bclXXs3mifgrm5gAL6mUhZ8hiVGC9oTwqSUZh9s/VkkCcqS8j9PaXY+VcXs6/4oCns
Uj6nnE4Owx0+fKXAds3yuYN6m2EUncm9uOsmW9ode2Y04hkJ2epJmwWYMTrRVdkCzIX0E1IAimyT
+kQzXxSAj5TN4FhVfNsUlhjxioltofGwEOTBXLzLkfzMMZDkZmamN0RAZ7eiuX3mMWh/RDalbuCv
1yupwQO4CS3OjT6hvAonuiWnQ/1Poqf8RsNNC1bSaf4PNH0i4ybNCvQuOpw7+xoDkMyQ+njTx3Mk
3c0PM4gAK5Ib/gLFy3L4DIPOaiMkpUmmFF0EI6JgXGZfoVxYSMXPc/vTNtc0eJBUmCS54Eu7J5Ha
n8UTl56DA3f+3a3eA4n4EGVZMDZqVYLfHChC20g98GLuha2MfA8t4ZJsPQcYugyXQWHcWlxmWdvT
t/7ruj3HUcYAHWgLEyViqC5fUj6txGLx0e2KVFTVWvz/mj5m1IzyLP3b2qDx94kU8s47DCHw+hqv
YFd0bjsbQ+q3z3WFMofx2jsw9+TFVa1+OUQ69NCuV2vvuMg5ovHVv9ERGLw8g+tNJ0P0wujG/0xP
qb2M+ov6R5/2NLSZnD/r53pBuOvoOyKo52SJGYXxOoGb4BX8xevK8Ge59RRaXIpY7sktPwoq93ZT
v/RsJFSucGj8Pf0avlshYX14CBd6ONQheViB0Wh5Lzd1M844HDx0XPxorXTWbNr07lRFMXoMFZre
UK8kVFIt1rFxVuZaMq6IChtTw9dw0eLrYssyWjw7vvh3Tibq6VlHTiGaIvMPTglRvgoahWR9D8LP
5kZm0SVkEqxuGoHM9ubDlHr0BPxYOxXU715sGU7JoqsG3kq+hJJkl9TVs7QjANTQLSpWZa2jxpEB
nkzgjjBmBqS650BJr1vRbjbEntqtGLbkaq9zUt0Wf8NiO0OXvGCBNQXyct9pbzGUvl5PqQ1jXhuw
OuWFkQhPTx/H64lMldV21SImwazGkCT1/Xo4GqsGzkG/V4zIBUk4+TytYzlnWKMhtvwXIRiGc3pf
u50kvTNIwwITiOtfnam30UTdR1sK+m4bLK3OSF87yWRZwaNRC+j+d6X1wpaiCt+Oa2hwkAvRx36r
7AW9I53NpcUpVA61HfRzTyAIqqwH0Gg/0j2qwW7A/4F1gFyXZtmKNdmBryRhc+tRVWtGxVjQLdIF
eNIR1g4ZKZ55dmvAQldvYDAwwOTD2rY5ti3I/XJ2L1S8mXTdzUt/oP6FUIjWz+1Z7wDd/NsH+qvA
gc7XQieZ1iACIzk2gGq6nz2NKolI/DfRf8wWVzKV0ce1GtSnY5Q3Or9JVHvQ5TY+5kGz076VbnoS
JsIgEsxgbCEKirO8Hle+j3+I/nbst06Igxzv05hBnf8gVrGpibsFLEsGGatO5HQRqCs7s6jVaFcr
0TkXRYAAfiGYdSoLiuLOnZxut5dDGd6yvL1ccZMheT0LyVyVtMyrJPyIaGDhehSbF4wZ08aYUEQ+
35zDBLiNjmLEKQr5GAcpxIltATPju0y7lfq+xSZQC8UsQgp4NjDOD7JNa2IevwBIYf1T9TYeRyRt
7bDYjD+ZMrL0lp3qxSKCeouv17lAa8aYysX8tLmjfZSvvA4Y0VsolHYOT8yNt+LuJVmdwv5VPztP
x+QtLC7+6Acw5kzftdcGPs/6s/KysK+mRCDkfKLDVFCFcf8/2FSC4wuDWYPNvyImO2Vked3S5Ny1
80MyRF8isEmCi2JPAt5IxZwAMDV6FsyBmr0EBiyr0Xn6RloLCi9dYiXglIbGWlZ70mfnCIrcQFmJ
9CU+Rc6arFbB/ZdfbkcVwkzgKCqkA6mShUiO14jlS+9AiEL23jhV8R3dJfErbVzKEyQ3L2RlwgZA
fM9vKs/qSCcWDBXDVtuZACNIwMtFEKneoBGXyozQY5a/at2/VAmvO1LjoHLCHpb9cugwA+OLE0XS
Fi/xqe+YinsJslBIM8rm0cGAHcGJThLaG6BSUfcT88YgelTW+BytptdgWZ5kNy4ImYxrHlfVjDiX
MUR+nMGJYuHlg7G0bbpW80KKjQ3Hplxj8IYGLQ+fnmXw9x0/XQKXXVoO5+h/5DWT219P5j1O1gPS
HzFEem0k6EtzAsMIq0KPfHpCYuZ3bZrhFBr0u2KxGvPGwX465F5WxiIYeUEiEAl3j1s1tL1fA+TV
Dwr2XkMvKpJO54FFvZiuQMCboR9NH4+NJ4O6B318lxRzbS6gVfeGLmabsaLUHQVESWhRDTxcRzeq
d+2syN8OezcXVgcgWkdGM00+hwgFVQVv66BsF9tOMSrXxaOmQHUf11s00jk765eQt+cd+fwjGp4M
paLtgKskZeOz9GBJtrjA928SmRUsh9Why13Zd4wrnMAnDUdDyvVsaQ6G/k5nZONHzxGkzNZH8BxF
b8fzYBSaTCFjgWCizR49ElTV2BDqAYqD+tcs9IyUpkS73R3rqjqr7XpEDcFxP09lrYiDEivitX5H
uG3blzqQKhYo6ybPpDQ6KR65K6OuOvIdIqrEgWeimNPoRXW+QYLWNildnXRqOfcf1RWhWXvp4zij
inZyV0TdBsYiFSXLXYegqf8CDjoQf6TrATugUd75T52DRmof0dxw4rNbXHpTwuj6WnigIA0HzjJq
xPtezaEsTIxvGq7plRxw1I1sOYonfkORdbJ2lpVgnKQYUqKdEE6oDkg2wSZYcPRUc1zdrO4hXTf/
C48T5n/XC7EK449Glc8BY/Qr2WeYUOG/XRuQsE77AUNyprOO3aUiFj0wc+/GTvNCyI2KRY3MQS4O
XUSJwrQNoTxj2VC41nN7dLxGEju0zttdnP7JN52Nx77g1Eh003y8Lfk/mSsaC8bafhx3/Xlwro3h
kWhaORbJ/WFCeOHFiTKrUNefh5lFUm3loECH8YoKpZiCobH+5kXCmM82LbI7F9OLxB98iwJSSBzF
2ZztQU5nPSRfkOT+QT/KD4vMELzGmuGJs80tyMocrfJOdGl7Y0Nzf/mL3B2+nCyVpx+QKEbGLa+o
mpkTExjFrZB/6EllijUtvlchcjTUvjOOWZFYHEE7u0CeHK0x9oyYgCi2qt62zTN9sW+nojQ4VHXV
limJ2XDB+AQF4puRpH9icgLMIglsPsdkDuQVEbXxpvXkWGOZHXBYJUwg2Beumwsn7du02ZeQtFw0
orCTfkw6myx4n3YMT1eod/f3Tx/TeKLqCV232/xTtnggODfaUIasQb1U3P7jecQgggG8G58hgiw2
jjJZuwDqeh98NYPso9Py6ylgrv7szEX6MPT6v4WDJyZgMCaPvBLZX+e4ukwq9jbOTIV/B9hbKTDu
Ms9xCrhTB2VgrBc1lzb/5bGc7fBNrGyRaG7kOzxH0CkAHbeeC+P6kWMTdH6Klw9yCvFghXwJ1Svk
c0HECcJ+PNV6ZPKoxNOtEUz7LezUBcXsKEd9QRw4L0lcsSCAThQG0AQSSJp7Sk20GXNDYJl5iyfP
dcy5VzN4R9BLqnnB2DEoHdy/lkfexqkrw27hV8anJI0GkLigTR84rOg2S+m/3TtiZNkK4oT4acnB
wB8KudiNlC4DRaIItxOaxlKijL/UueNzHbjEDzTNrJOKcUtUvSgTX7wE62aWtKdMPHC5x7bf9anz
71+DkzEUZPLuslwqsY0yWAlHfSX3fw05QSmDsbaOcRc7rGSYw3GX7McPphmP+Q3BrTD3CklRKicy
PQbG26Tr7XsfcsjwrTRp3ziwN3Jid7zulqY9e/4tTerGce2ob4KSBnJsxLTOCNZY5+uR0Bw2IaSk
PrC4IXL5h6fdg6im//pCBdFIoJ/jCAXNsoZ49Lv2NNjRyWhS948d3VFVqLSSnVODwpa5LTzRrXMo
nWSBA8ozidsKxFNCRaCsIZmZbxBvV5vIvdJsFWprR6bzycZmH8EvlfVH75+09IMP7gBOsl/FTg6K
VDKjDQCI/AIymDcxS6hQZbutlF47/ql0itubiLxSXLReExxkfhJq4nPuN6wCUMkc2lc+PosD5xyL
LswGrKLqkJxZ49yScoti8KuOXBHWLDXDtmYynujwT03oN9V7jHY5FO1hj1G5YoMVIJMp1CDQmrcf
rLVvAjAQnhD6POexNCZtFwmlUwYmLKTUvZw226wGzNJh/55KPYqjuFAxv2oQlNnaMGbhcc0jrF4A
r7Aax68cZbzG3ZIh3hAVwEPTX/EjwpXrun0zhPk6yJnz6WtWlw0UuMsYk+KJn0LxXg94hgcBve8K
3m87AasVR2kdb1c4bmFkdaawa7GEQ/WhuPzRTwcWEKoquB1MhmtXXxEVSThCZ20ZyVyNGtUsQVv/
YTDthTFe0sj72fGussClzjcsCBPw+xZeDUQ42sR76+RmJ39nnCTtlfsxqxCSoLVb80GYCP+e+T+3
HwloOfZPJ/3Awfu3tje5QUrTzRkPgcxkGDVOJQZdC+1c3vSCDMpVY41cEfeGRZqRzxa9NgjI5qUw
ECXjjs+bT7KoE0v+K85K4Rwi/tt/g84uF17KHrVpLavT/N2fz8FUcL35xHLvz8c8HATr+sdR1zTH
vHe4o5R1oyhlGsTRS+MSWQ7nj2E5lhl3l3JkkB/c/T3sD7dST6zL01tZkPHHawjs8v3pSCGefHTc
Sf0hGsxku8H59fzaxkh6ZfHTYe0HhMqZKvUabLz66aAiuen87fFPmjZX+VwKT59X4qyA5pEjuwz4
P+aRLOoRlyhr9Ahb/FtuSa34hwEYCOri7H2cgDqx7MQLtk512z8J3rkyhPjqD7c3ufTdr7BaHpwa
NBnyU2lnyF0N1lgZb9axKDFKhwMvh+VNMC4LKMLjnhuC0AwIFws00qVprAS4kKksVgMRZNlDCVN/
2mk6jPKzLNnHdzGzEWw+2REFPD5nhPu45MIaS7y0lqagCTjjJW7A0tKtQiXcDqBPRw0/jjqsxQu4
MB1fNyQ1hvNHrf9TkXAD6CyXfsNqWpay5uT+Xd1EmID7j1bAGY+qn/+FK3LvYaWLni47gH38znIJ
1zv+8UbqG4A91u9SugAHNgSL5iq8VbrZC2eBdSqiGhGtCvnWRpXrw2OZfWO/huzYTs5Omdke6o1k
NWHDmQTnthyRxHDAdIBqxizo5fRe+1r2EB4SsBJjPfQPAEnQmIehhbd2k0cUPkMYFxdjgx2YUhGT
nrMKTiY4TE3zVBW+FOuEHj6yhS3OFgpudK6R6uQpt/6WQWNv9lIt23hwqyi+aXr/1Iwp/bkfEPRc
0lQ00Iwb8MmhdiJfa6gxfEx33EV3v0wdvb+IFeafo1SHGU10mnPMuhl35AFRN1AsoRkvC8GumQm8
kUv/gIJZgWL7lN3t5Ortc2hTBhCcjfQPW3JZTooCj1PO5gxAJpCoefatlGo2JVxV+i0AmKk+nMXG
04DToenNCY/PQ/PQU8vDNilQYWXr4Pimu2lM8j1ymyWjeJBlZVNP60JOC2INZHzcaugVegjYdbUc
JS45lotoCnU1RkjM3GCaPuSbkQPBxn2MDZhhvWVUlMH0MTi1SkV7gdGwpe+XMKm2LUv6Ee/kQ1T4
YzVu2tD51MaB00wMtCiE56oiwjYxst78FFeAoIkBx0TvX1ylP4vScLK6al32jkm4CHciVDiJiXIX
5Y+Maxnrwh+R+rW79MkyvI/Fmqwrw6strX0UhwY3kxK5h2DcMEDYCpKDP94mTEJ66H/548UT8V3n
+AyTCdQ1MC41e+QONhk9hQziFA2FNKDH8an4T/Q//PnXACnuQwmGy05/84mexnGEqywylGCZA+2n
7xuV+0TxMYw7VNZjx4JamaQRnK5ImgQQdy3PgUfLpofJ7nzp6Fk3vKM+e40MvnjuX47a7rsLmn/q
hD2XscPzfoum+tIadrJOCu/8n1sY4R8pezVnKxRazN+PG3Sxt1AO/XV2Bb54Hw2mojiscQ1vdUtk
dhJhaQBlMfK/GfzGaGOkdaeGw0m1eygE2BrYW0BU7DfynCF806XprC3bMeiBD1QIWZMLVc0jva0/
49ZB22qqN6owzFZNcI/84UG28LRquccORmznaBNV1M6hn+8LMV5+ZIBOohdGRK0Bj/U8ATHBXDvM
460Jp+jU4qV3CxxsAhWXR/g4IVky+BazFpZb966g6lEf7RERs2RvtfC3HvJ2gkJj7X+yN8IpafZL
ahaJohUIayvabBf6NKRpGmowomLIPy60YES9+7G8bJQ1R0x7YosnQwf+NDvSSQMg+mzMOtUmMEJh
MExDZxTt2tEEkImMMiOgq5GpxF1wh7xdcp7n4WyfRPbFUnQ8BiIMnIqo/fSSrqqm/X64GEkzF1c5
yH7i/DZxfMMeQYMqO5c7iw3EVVLzsPNb6FFLpffJj0A5tyqjNVLH6DjnC4IBze7aZ5memkCEn0jc
c51DqetEVs1HUOmtbVo+hWHQTfgnT1tbFFhVQ5NlgYxxLKXGBfXLpDDWY8u7Uh/ts3dMjClxj/b+
vOA+LEPWSb+UFC+T0qOXFXivbwa/xsOQLv2KpG4aPUAEnF5RVd/V9VqB/G3ENtNmFu4hwu8mB0f2
BTnl6aATQLN5SbPKWCV7SRHtngO5i/ZzWGdCI65TnnvQM+L3Etsq4kmgMoCuOpmC4M5Ldr9h1YZZ
GfCl3tjW2Zn4+jb3XHmF8R64VLZB6JcZ1VKOyWpln8tQ9mlSjYfLRN24/PkrskCTjcZtGqdK2ZOu
Trz+RIzvk2ieV+GVVi2O0PboPPpq8Nk38+RH7KK/kkv7CPSSnZ1Kkd1oEn8QWkQhtgMYYqWGroVi
uwvJqGW3Xaw9FgmMIBFxTsC1qextTNEN8kWdDbc7tQ4D95cBEbyrysaOWQ/WFTrY5nTDXWn5Di8g
5eRBfCk//HXVVk01N22XVJw7FqUlk88ARFKpSTOt7FsqN8ZHJWqijsYhtc9nasWatrtm8rdxxw2Z
5ycWhUxfNwzkKDvw26la5/HOX1fFCjiqdz0JbC/LQUf4LEGt6SZGx1d1rOq3+RnFAdnjZIdnyKk1
zoljTZ0JP0y1twSuPeYjCjPaS36/l0+a27M1Cd4+q2uGpcHl+YuXGgebD3uYO9T0Urqva+fk8NIf
TaaaWRppObX6uDO4lSg9Th0rEH8+8mhy3oFSTmgrSorXdmzbCsS9OJuSHjYMae3uOugZNTeW6er4
mo7pvakRgDmc77Be3KplMev9x1++UUBC+10ZOUzRiH/Ufo0NILFJCyFiRjNX3Wy+iFwiMxVWhwft
ow7J5Wvve6Oh4QZrLKddRWT+6ck9oAL3dyyeM1mjNkSEidE6P+zHqGIEdNiyA1X3ZXFxRgAxhb+L
TCSiNAmCYj1jZ6i0grNGzmnpdEOCWgD7PDRx0MG15uU5nvlxBD66FX9/WKFxIoUk8sxLYErHrzQY
FvoWsuspPSz0xJxzeSPGOYqrJH2tvM2dWsfWPBB00rwDS6pQnwCdqkKI6gZsOrHuu6sW/1Asamcr
uRHUQpN5nLKVNDW53VWm4JTD1YOVWGlsnIVDLAKqpdGPh3tTR5TR/aOGqBbDfmebvgUzm2l40Ojv
2CmYx5mK82g1F4RPeI0kIcAun0pHj2PvnLSgfTyLqNLd1nVFSObr6UkSluGEE9cglDfavFRlkqlW
BjN0cFrLO0KyOKOg8rsZHHI8TnJ6t2zBSibxQDd6q/5R5kzvgT5MNgEQ/Ig30tXYvY7fuWpD/mtP
mU/3JUPlA+ReeSVACQmEez9EkfMPh5T8JbSDTjIFKnh66vDh/P3i53uSZyPP02vDHpdW2WP0zy75
Xvx6bDzrNSpwFINNI+SMtoC1fwhGsA+6AKN2UlZ8xjpK1iN+451FUqfWJGpc1wMlKeXgj/djyMbz
lB8LZ062ktv85DYFDnXoWNXOEPb33OnU/r9qTnC2MLn4Ynks9WAHxxX0dQGrtSKOjISTuz+EPaDj
wqsI48OsD6lqiZ1vw8W5hzh3/rEsNs7aQeVRzlG0kdH2x1P9VFxO/uZe0v+0cW7GkIii7bl+z87G
MwCBXBvshAfzPmuAwg4+EMYRWy02fhYbKgx4b/7LQj69biWv1tVVESfIkI73XJoqf1Zxh9jm5jbS
PrxRoLKITiz+fHrFH/0zDusOU3ia/LC1tdRwzkR7UfyB5E/VAqvJq09zCg2pJObBgRuJoQi9VsXd
DX1n2I0citsVySzR52N16FCKtaNoBJSPAF40vIyevSUezNC6x8a90l/128P/MVdNQf6MTPSw9t8b
sMUJqz+ofZVcL2FI6wtlXx3hHQsQkHPTJltq31Pa+iu41BASNfYY7OEJ1mk5dGyEvo5IvzR4RYKf
VszTu9Uc0eJLWxWshfB5cOkq0OuNdY8AZ7y5K+ZJc7pCGNPeRgFMjT/sVXT5rtvKO2ttDi/sitUM
og6nOEurxPyP7og0E1Cd7LQyNYmirEWThhm4Z4lNvQFuQEALObSGq7ZJ+CV/YWy2stUw6mD4BMC2
Xa31skQCdF+yuMzXsGrfm/an4pVbpcfw1BHf63zvBhJW5X4Oh9VlVweEYw+KzNZmmCvgnySKLWoO
w+1Lb37TgpZDa0y+UVyVrdKOjMyI/QdQQL9PjciTqPmWk3+okGfE6weSgtPg6wuB3L4qeCrOvhIb
gghHFfZw7NmirsHkNI9d/FRzk6y4qd8lEmdsAlkXZfbJbcwihMJLBWp4qzAkANt7hUnKByFO/B22
HHpGEV97FWOGPUTr0+iYaLzDHqhnM+nhiDrsj/ofwFVW8DeaIJ2Y+4GAlKSNMz3kokJkVOV/zPd6
hpREewEuXM6fownYYon/6gxPDYVm78Gt2ZvOqGBdkJ2GmuTots8fps9aMjpjQwVCaM5rTtzYGP9T
3lEm+vScN6Bf9mZ8h/pREqHk/Nyu60JYewrCw3muW58pYCQHEbyW2kZ7Vgv+Jj2ceSM4Nqo3a3X0
1Rfr96VJ81WUvVLlxZoVUCaT8yjS7FwNr2oYgb0Dqzr+5u9Gz9gQiOwUsLynQp6KU7rbIjaF7KE1
kdJz9JZ69yanm6QwhkjRk7B7e42urPkasFTYKRXhLek1bQmKnz1DzncNqtnyOIIBdmuqribz6Ujb
hKpfsSBUO5AIp0QTr0lhK8uNTprOQThpsA7qMxCsU6IsNTFetylOF0+zIAkdXe8WayUhj0i/lKkp
uAa/QrR08cTyoCJMz19VCMo1E3EMbnLN+u9YEiQKmXpbUeO/GnkbKEskdmN/FRbyhzpA/MjSb18D
e4+U+ZR4zeik4E4rxqZdVZ4MCzEDfXXN0xcQHOLVOMtGNMt2cFJdsdHyZdzL6Da61o8aLZiGXRdi
FL7iU07G3z0QF2M739hS+c5gigQA/4GewRpHWis55ZSesa53TaurtjKo79Eqb6XZ1VrnYLcfYK/u
ZpAxTQ5j/ucq0b52FIAQ1qhKsSt4PqGhjoJSIFmYdEyIzf1xjMUe0GtfSX/nF/X9L2/YDPHY3RDE
BIakNOTl3SxiQ/L5AcuXfsXQsTo/ByLqzI+S1qhf7Y2mAOCqXkJwYXBEBf3K9V6bgKuS6dAE3IvF
Tm6r1GawSgQnEdX6SEOUe/oiJkycXLGLk+vjE5wW2wZ/Hk9/OhCK9Xhc6zkWhWX8AV7nu9zvbzne
EwLaR2PPvi1thzgkR7Q3rWWwYC1LzmgwtMxc9dkTXQPXFIE1exfHan5h+nyX6ktgVPAF3r4zKM4X
KnZQSiC8kgW/sqtgkKyMdIXizY2mRbYoTedqqgMdVmHL2n6bXhhQ/bPAMSkNXMalQ2dbPc4uU0re
Gb75vFs86KM0y+QrInG9db/ej1qt8zPsqJPN6kEeUrRjlLvyIvAS9rB9iWxSVrbUMkYeHMm6pMDP
lnxlCH61/FdZ7x+sZSlKNa0I1y/OfiHIwDYP+n/mYXe5VYr3TSPKdBpruaUiDUc5v44p3zwIB7fc
W2dLve66h+TSLGgM+fesyheJ6Mj/pmsjY7YS8Inpam3vE3lfLrDjeFLqgOuojZxsHmC5+isJbH3N
DNUysxQ9pfgmZzRk0UVXcdTBTAcnUQ8o1sKYbvsn+Eb8MLC0nJsV8nF+WRbX3pFnlmxRXI6iXxq+
4yC1Vq6GJQFSML6rzlP8xAAOYDCSxZZSOYVnsSmM9IUH0mZ0aq9Wzp+ElIuS3MnYFAKElQZ6abYf
7fXFyXDoCAgLGHwkBQ0TGTq5ZZr80w+zdrWv2+9Sf4Dl0pCBsJerCPzgNgk7/oKSVitgAJjD8R5b
67IpjGLiGP7FN16//xpda71yqFd1FbSnQOAcKZrsrjSCB0ol/QJrVZ0zoXWK5t52QC7rhAbjbPJx
1kxpi66YjYJen+yao1DqZMY2Fwrt1PUMm2J+luJGlr5QQyjjli2DHhY6UsFp8EoOAquOvim/SLkK
TSqAhAZL6aTVX4Oum7cbVcZucQLBtrDkn1WILDCkim0EWOIOr0U1fehPYn96jAYwLE5mIqLWblIw
Lj/a5sWOrGEuue8gGBv3qBxIjficH0nI/+RqCmRe7pU3FCz5E5LdlvzJnnrumSJsH60Wd35239j4
Bwdk4C/jmJIwQqFDIlVH/2oTrqTDVCloRWb0NO7ZwRLRoCJV69lJ2uVASdcEm2V234mryBrXgGYC
59BvPevaIZnqOvJFkqld444EHO8rBGwBqccK9Sj6CCBhJgAQf9rTeWv1ypUB3CLaLIX//XK8nPhV
h3MfNh8VwgXaJnJBNdg4YfUm79YKuOv/oG3/TaHJoTR4c5w+yYscn/Jy20AqsHZkRWnCCn2S+CGS
w3Ks/eGKY62vhzhCMC8plWElNAOoWb/BALwy9T061lChjGRUBSuGzGezfV1lGWccqHODYeysCZ6X
9pk6HTsrk/OI2HgbvxNlmX8pTwbd7/911YvTluvogz217rxPuR0pVsB+QwFVKnf0ItcZb0LMX4uS
plvS0pwnG8Q698FLv1tIOS3/40H+fmbGH2P2cSkde7tMb4Bd5wkDOHapKiOkxmM0ML7y4FA7v9ND
Pg8mddqzMap8UQA7ATz2diDOcgZ0HhX4/o+jyGwKEaFRgSj/yT1Qzv7EX9cjM0C9KYpJ6NofEOSa
XFJxcP3YyuIPvzeo1kjdpv8lx5vOL9bmwOHDXRMzt71PXhjwMOpBWYzTXhl2wyzrw1jnyUufWul6
6Gik9DgtalPJFLs3NrK/HsjonkhIv910VIeDqCO7BHRCeTeqmHke2C7ahkoLLRazCT3AAynTH+8t
4bleRkxKoIagrKM1k48xd/T1A5YpfWQ8UuLCiYkBbAceg/41B3VEjIcj2rrYrmbRs0d4lheqOiPl
+bWZg3xmIptNMwVUTGMJCHPjNhDvhx1LSFPjKvnyoBSqM11w4kUYHYBYnjWrg7M+vg7NzXbIhCx+
F/qyYdc63Bqo9wl8rNlOra34DwbBCskoznMM4HA/mHNECxaowm9abgHaSK67t8ZoS/n5QRLdpSDw
o0UpRK7hA/TB4GE/tMxZG76iVEe6rNlSA69raN1i2NvvMrYwHU6h3sVCTfwk7ozlh8Ar/5g07iRS
lkX2Z4behlsUJfB6wFmEpSnx7+U69R6ryFSXFcn5sZTvse0mRi9hQto8EFuBYrtHacuy1VkhJZ9q
3OamMzGOInFWyrbzkpK5OZhb/NW9bIbUrscmOmuMvXoP6Xc9WdGRcLMPFr+O7kwrMptXQBcadlg7
LzWilmuhABK2kXzRmw6dlG/T4kzq4C4NHzGtUkM60Usm3sg9FQPhyYTuDNSFM379eFxcuOmzdNnc
8gdq67S03cUdRNkTJDdlLWV1KyDg2zezyvRezwKAbGC5M7Lhbo582IF6pyod2guNhEzYK49nfoAh
vgXHZXDpx5diE7FuccPnozCnf3xHGqNVXGGcx/a9aJNWxdBk5BLzJ8fsqfzQ/8SsOYQhU5VlDy0C
4lUNZRfgU7Difv+UbEfFdaJNrOXBDulv83YmWmCoTu21c0cq3W7sLLCCDcvbvqN07A7mfywpT99o
ADbFBCrGMGfgb0PksTvZPuCzkIAYaUlxf3MPLuDw8dzmsA7bYjbroubuqaV0bSlu48jXjHXxAPLe
hcAbXQjbvZjKu7QsOcEmorbl21m6uCyHSHOOZ+OnUOcga0BS3cb3izBdFsdXMzEN1dgs4oUFhg6/
ySPAfZsCZy72Sh1r/jZdHu+yTu7/LtEIkh+6ri1qMlc0HBLM4gEBr322/7axt+zSOmW/jCZXRhS0
W5xnMpNJdrpnBHX+fxl7BhyEE/CVHvqI6WxoDCZ5zETuWn8Q44O+ofbGrvl1Nh1G2DlQvQJ5FE3t
sTFHxaltKS+yxV9bVij0i6L7RmmQ2pLjJTj+nNRMWJGByvps9QuFyD3aqSe3RKQMuELWF2FV93wG
dMWrLqRBSNpWp0qJi/sA1Ny0C6VGmVDjZ0sQz4TMwo58dKwl5zxewiRWObE9EvgTB17ksExj/Vvx
bma1Sm0gY8FgA41OIGFGo2BN9o2u+oda1HyktnUqYFCuTl6jW9i6V9ioQjOUbX9geKw8HFy8aV9H
XvP89L+Wyzm6zETUlymqCCFyrMNgxES1ODw1Skwyqia/6hNoyW2vevAxnFaeVwDKfH+oWV5pDcMY
J87GHuPW4pPFELsXSAs3/taEeyQfq6UsVAXLFGgaFDcKKL0JVBhJi0kdF+NJAv8aLDc7pwh5/8yE
yVP+L9VOOtZwTaRePIl61rw4xQ07RNhy1rhTCe7gLuskTcK/NQev8B5p/RVvZ7+QBW2imlkizNzP
Ar+3CoDFxxkfb9/puxxmOrmo7seRVmyLWcpxAwriPxvGXisSM836KGBcDhv1S7635U/2G5e7w64o
sAKnPTIHMO7lfZrkFpDUD/b4M5zXovs87x0Jkqdv/wHj9wLTIU+wrvggR8rPxKz7iAvCg2DN8RVd
e4Hh/4TDF59QYe8zzJmF9WrzY5que5ncPWDjrz/GihGRNsyuxM4cca4qwQP+94yKllEPJflA0wLA
AcZ2YyPwJKGsd6qk9UZ8ruOV7JY85mEOzu47qWF4QdUwuMUJOAsqsX3sIkzJ49SC4ElooMSeUQ8b
UhOCPn1cpHOExz/7R6BgTR6GbRrlQjC1zD+zDRbDHqKp746GCfnaezNIh0rX3Bj6IxscA4P5KLAE
69c3XoA0fbxVWy8iipksCuayzcoRZPhH+U39l/PdUd+T2oiPce1tPNQbXayYSEetMmfULl7qkpJm
Y64oGuc3Xzz/+DvhRYl0VF2Oe2p4Dfvhd2TRBY7ZphIznt3xW4fR23S0jbyoS64Sc3C0yyUku4nf
SFIuKxpY7ilbwwwRQIFlzPQVeDrBryQ6ceLmWAcJoDhz7OEh02cR80Bd0yuY3h7hiVy9hXAfgh7W
zXOuxFNLAIdLe6ouuBSVPsa89rMN7WZFKAXBmfJz1eAmneEoh6DdguQhNB//WeHzFE0UQg96NbjJ
ChFNa220jLaNJiOrK3HPK/rQRcZQK5lIIs0hnZEpPG8n20zZzcwJZLq+WuE4A1liEN1Uyx1ZrhNo
UZYWQ/KH9cQYM8BXqdW8nhkHzwhz/gHk9q7YyOronIdSrhD/RGsTQ1gaL/sg+vSMC5JLRv5N6wyx
EHB9FoC8+nKgJDTidAZ2D29mGFrVyzTAUTqgvtiLDTJJge+e/KIRrV+tgqfwWC+FkxJ2LvIBKAur
WLiDM0felOJGJM9+UNCaPgKDaya1T3wFcKcBlxqJ2dxeQX3rOe+NdvCpRm1q7JF0EiKFkniE4lCM
8SzrZaCKs4XNy/u+7q2APtCedSzdvgTSqtNEEh0lIWzFFUgtD9rG3coBDJepIDff/pVguOHJYVE9
9heA84hGiYJeMLULRjYMcA8fEyCc9z3qFMeItFvvD7ZvrjTIjbqDDjYyn2d1tXOaRqh8jkZP5Wa1
h5WTtov8C04NA9KQdfBkhrVOKv6s79gqVqcygiNnOj+uqBdDdIzPTLn7g/4XK5fHBiEGuwNuY4QW
uTdVOvfSoHkta8/Vkhivh3UrnnNynwTxmyTXVHrfHRNpI2JXU41VPBaCFD7dSbgC9RcxW5Hbgej+
ffdKWPYtBmDKKo1VMSBhTIbNtGXiWLEwEBoxyZwyPC+W/EdfGvh5qc1ya8G1VgC6V/dS5vWyYyOP
DlNz8vsjuVVkZP1TNNAHrEfUkLoqh5yZoUQQPyb84JGJtk/U7oac9co0WbdE2waopbhtg5yQeW4+
zx3d7i7FiQkyA54hsCy3xwDKVFgHMj5X8EV8YE6kW7+QWU+0KECYj9LzbNfIlnPeZr9DO+UQnCxr
RAEAqZg+2SKPuCsgn/ofOwVtaqLCLzAMaTMP5mi+TSsS72548zvNNDM8K9sZeB7+raQ67rCeH/Gt
kDTFAW/WnHYAr6qUbx7jabhX3MRcjVgEEHCyUF1vA/zcNr5AZEmEugySyJUPZ6y98QZAcIDNuJdL
F4YSrLMc1VEjFiwhWKNPY0oG1glMTxXz3PFrydFNedfn7ncxR8Lm1b9qnYCaOfhLR2chhbXFzntK
4vZihVmo8zuwL7xJbjCc6DGlqPQkWySK2iuUvqS7bxlS0rnPlg0ikrh9dw+SpwZMBWXEDxDwIiw5
+wa0LWb+P3vJpacaXxqb49d9PyWCm+zRF4EaKQYOSvGgLp+Fxs9ClSgPN1q6d8we2WptssKYbzyV
rOFMquH93Kn6SXMx9Hb8bwEVpvPsQlPcFtBT79w7bJOkKC9R21S0uOT/4RlmKDyvBzMOJcL6Y2/k
9kVBWz7uCzM8RM6gw4kB5Q8ltavmv3hnPwLjqIw5YIcsm3wK4tvJzIvFpbYB7Y+WUkLkTmINTzA3
IuszUc2kvjHlOunE8mAU8HFcRMx5MikG0OfRMQxlzGit0SiOHw9Xe6K9nW78DV0gjsMaUDePMCC3
6t9RKXS3LMgPPiqkf+/MqRUWIIfWsZp5nUfUtwh1h/f743SRD32cOyst21EFm+fgwmZRambJZxLy
UfE6j+mK+RqQjh1UZ/4JMAcrqU3aq0kaw2fPuNHZF5kWWhvmYCSppqDQK41L1o+vGpMOKVyU99zT
mDofzciSu2ozSm7MueDWvE/vUmqUUQ1CU/+lmveqxl2c+ByQjWP6iMPOBsj6M1nI5xZe+buF9Hls
HkffNyMDhSggsZmZ6YDZi4mAUiB8hoU8p4IGaXGmig+TzLejaUAcg6Hpv5xISZuH1V8sgzCn6OWy
OnwZqKXOIAhVE8+sRYT/DpDmdrNkl1TxOeZGFm+tFIo8swgOCWvupWx4p2ZC3gvyJs17YXNHy27U
aflktDBVDf8+iqHjS6N9ECZlq2R9MzQBf/MN1t+FiR4Oz36t9X/IBl07/w4rybR6WdCKFIoQBGZu
cus6ID4ncvRIXyRO1PQmXCIES9SnUSil3wTt3awckPNImALf5F0eSK7zBcmdaS+uwER09WEGeNyp
fvLOITLWWqyyABA0yictwSP3YTV0ftEtQF3jOMWTzC3ZdcSloXRIeFXroAFlpjjqKFlNYu910kMn
B4S20dYegPsQWVIYnCwEcne1pBuPBl0iMGM0oZL6qsGOGl56s+Jlv8pqD0T4JgyLTaP20nwUEHEc
GwXDsXHYonV/UiXJ4WJLlLuQlcyZeLgJblzEC1DM7MWCPDi2rjKAFm13ru5sDq8RcOlUGsgUtzJU
sNpzSWzV5ptylTfrego6t5Zif4pGhyj/I29QdeId3GX/L2oF8pOcbiOKUdJlFitKUEkrlV3jHvlV
fzyxvc1zeS23KoOu5fdchktlq5dPPHF3X5i4TaiRVkiJy6FhGevKjNPCDkf/8om2qWPIhrYYmnwc
h3BCmZOcfPLTScxRKGf9zjaBP44paz+5u2ASc1C5XaPAnoblI6kZ/d0HxOo4yBWmey7EiofLifkZ
OH8vdbK45+zBIjvVkUtxSu67GMZTtcVCe9qthQwDfys8KqEt3v7TXCWIrPDFIaO19lj/TN/7sx8H
2xI+1LzmuCtz4WPUUCg9r4CQ7aGxbB9EOtKdoRDok3AdhO2ZzJTWDCy7CSK1qpIAhrdQtjhYASkC
DivfAdZ4Ya2dOO1fZvyZtpAOzY7l+muQuSMKJcxAqfk6PqYBmnsHsuJwllcucexMWchkSXLYhylf
PSerK+33CacgrxsvfoJbohtcIHgcdfXUdVYHeU10Mp8ZwPiBitABTJOKEX4ZEXG0idEScYXnFDXV
jX9FNhjbSB0PWyD1H/gReAV+nXbVl1U6CCzbK51m2jbwYKTOiN+U2766uyTpmB9ekyqgs9DXHmqz
cBLT8Azq9svrQ1XxG6udL3hcKf8jbYCov7SHMAvv3XvsGAG8LtKCnFf1F6VYLPxr7LgiUc8P0u1E
irc5Wy5a5bh5cNqGqAKU0vGYPnB9cDodTo9qWdsp+qYL35q5yKnl6/rkymoxkusl94YkisLdvPoZ
sC8FSIeVLrpy5McE9aLe1wqlTyzAN0xtInnSwMVwi2KD02EnOFb62q1ctKDgE5wiNxjfpq7Tbmbm
wZys7F9bh88DKCJ9Zj2ZYlnmti8Ge2cTBHYTgUDREEmyzQdoahdcV4vaeVIY0N5tD2/5rwiwD7pT
CpB4WbGYPIneYHX16B/UaPr0QZtNqAhxEnz1EC3wXNhK1XzAptCFCkDNngSIGCv01Woly3wHTi8w
ZR3Z5S6iZ0T+CNTECJ1I+AO2UeuuyamOS6gidTLQivYpHMV3Rn5djy0f41scETjiIOOdHyErrY0x
kdgU30Hp/3bTo2HPOh6EtDMFqxwRyRe4xAn0gHyzQZ2BMsYhrbvEGyoU39IGRBtSixKQWsPmbAr7
T9VYaMjcwhX6hLRuHqXJljpnxPHfvE9Las/CLlORlRVaSap6RMagdPXuV1dTrmP/3VqSiJA9ZHBS
+PjxqCemrQ/DQbDztzD3WxBKXG+gF0vC2nfdBwXwBg9MBTl9USDq+/hS/cH1KeV7Ep7MvuKYkYXq
g4Xd+9TXuK9VV1SMXYheu0B8xTKoqVcDMfCQoPY3j9hab90Gm1bqA+Hbfi6qeIAqjDL3msyDkyNz
WsSnOcZeDtanTUNMbe2b6aR97RDGJwQppBrF4ABLTOJbccvGe6Jc5AS1WKGhZn/xHd45++oaM6O/
W8rw8vbPSbHRkdLs/chWklu2nI2oaNq3XvhNPoHt6PEEQhp1xoqMpN7kovYvYHJ/vpovce0VyeMB
51PpSM+SBnW7zLsoBxGQsiJW91j1HS/w4letikTktITOJNRSoF0l+NhD3hq+QsQVgWXoFsV/IjNm
MC2zH21cpQBZ3e72tiKj57ATEaju7l/HyllWwj7DnwePmRjjPSHzK7cUQJZ8Rd1/vlcwg7ckrV9B
VKdQNAktItlT5+sfUF5Q4Y9AnfSUVieOwZXDjTeXkNOKy3EGgKwTUxb0/eL4rM+VJydL9YGgp4bB
g+6O8RG7lu2lN1sVQ+WIxBUu9l0aCEkAlDaMhhJMawrkF9lt+dRzvy7Qoitwymy59VbsuEd4bBpH
omxD+QV/zwBYiC8Gt+7x6YL+S1W6GvRpMzz8Dkv9DSdkdQDwLy0n3FBGuIE0H7Sd7ylGj+M3RdwM
LfLBFrZcTE9lQt4nXoIlFD1Qw3B1CYVEa7lo+gP6d6Fbg9DRfHviF1yTLYN91sFP61bQZoUPlf+O
TINk2HduohSnF9SbeJgcR4x7J+gPvd/uBn7/6PqzYnR3ll9L4vW5ejnIfZ5QugDy5S7vsr6Csz89
arIpmGCFnWogUIdqVfN447qi3/1RIubx9r+ywuA3HNb3WOo9W8UCdFLO6kO1PKRVNvEwpOqCp+GT
zcwMtyJVQqR80WVmxqIgmWT26xYDan4R0qhe3XceKe4vv5Q41+E7f0OwNQmrGfB+eDSz54MLIJDs
PYkNdwK/x3zpeEjreh0WK1JLqE+jtp1yCxEM23CRkyI+IojBd4gyOmFyrUj0okrD6dNwNxVqfD3F
w/KlpvX2O/PBmzL4n5gG4eP5zpdvQCoiWXX0hW+QdrlrK/33v5ZE9mqdS2R8TtRMSb/Sy5NZWoyq
+WX8G8/1K2zOdgypFQXqALDO2lHIewuPPyNpWHIN77oBTTUdBK+k+3V/Ut2R4N+idjBAQU7ABMkH
5qJrMN+bdKk0nwpejErCTs6YdjsO5uP5xyaNd30n1AnwO4AYtZwNzjzMsywH7/1fuzmnyP0wWStD
TqxjX7VGBva2Asy4lplmQSSsfBkC/hjo8Tj0K324BntGt3QDZb9kR+iLIO19gfDuelkANixbLwDQ
McpW+x5n7/DPbjOW2RBFGDnt+o6ImT7fIskX7jzWgS7bZRNC2k0NCyQjMO9FoVJ5GQOUdxFy7D8D
AWzP0io0X64FxldLZ9jxGksL0F4pmHEguBDr7OcA3zbJcqjNTGUb7458sKy8VeaRCfWVMDDje4RE
G8CKMgoZQLJ4NlLglgsYpl85RDfnsJaJRrpV+T/YvLqBCcjcBblyT6e/P6GqvBUe8vg/mPqRBhg6
tiFxEnKGshmPBhOSqphn3T15OToP6B7IC3MtWnVG/hii5YRn4omFnT/1JAKuhL2o6ezxE4/ddCUL
s1qOGg+YQXuxm3Rq2voUT4qlSdEu6Li/wXltbdGDavookIkMUZ7YmYCg1vF2uOTTIs5HphVv74B/
B1upkmQRUhInIgzDZRdYsBIzdFrTWocycvnqhYPWX1/8FIzNTNpb3jqd7OeGbN6lY9f8wzbt0Cov
GekIpG6XTFUZ4FJWPxv5OguUbkzpG6X0D1ls58lqgesfupCI3QYV+NKUhBgbhPhFQ7LPAsMExt43
NZ8srOGUu2pVuX1GwpDw6h7PE38xB6acTY6l261plbOV1YrKlKfV6z9oIBEKh6rPWLPCGTZbdRcB
padF1aWv9gW/YdGFcmFlC+l1oEICsb9o5+yRqC7D3pVrOS0y5RT1ajMeGGmFcMTTdlcp30AbVkNw
DLju+qBNTOG4wbA9W+8Y4t73qLBVW8xrui8Gjzom1yFlkhwky2zqtFSHOI67Z4adIonq3gTtDTbS
T3woUoH3WerhVLRF6Krtv6JrzrAumzHdvOEKoN1TLT97OZSrjsEmC/9R5IJyPTxm3VTuOIFX5X++
aMXwR/zee0/GdwZ+vz3LurviSf/4Zn7lQSpiyLiDMJxIOywkDmEueeyTWFCVM2edLY8tS4QsoJQc
Z3X3IEtyc/T1//MSPGDp4/WOfnKgezdD+kPxbB9xXUv/j/qEwAw1cFi6P74Ekxhuva84q/jlbUIK
CiJm9Ksk88e/0Yf/0JpkpBfPvylu69wXMUw85IYgHWcAsxDXWrHgE3vvh/QMBnZ9kfq/ip596mMF
4uumX4R54gE6gMRgOLP9B+cdLtFRFh+CjeunbRqHsSHF7LKK44b+XQfOXuXKioYuQwaREhKOX6jo
zUCL7wBSiY2PCAHtU1N8TwQ3YKfjhhDbjYmAuUEDlcjKgpyIgXFmnJmTZATmmFK4f2e+sShTD72u
vNS+2GMVa3LrJSRJBWgwEDCm1bB0b8miW/dRdbtuWDLLmv6VW1gtjApPp5YKkBGCo8yiOauNrnfN
WaC5GKgpZykr6iuqNNO6NmLs7Lc5yR/YJYDII61UhH27TYBAQlh9KZPhpB9AEaowJ4YKZAsukr6a
mOZfvgyHjJX+/xNiG+yf0AtI2QxaO1ZtXVh/vTOn8Du4vmD1bRWtCIusAZc4YzmTlbt/7yyFCx3D
bNJdwNVRbvYQRWXMymPsdG39VtygUL+kJ2MeQKb4kzfAawIWTSbi1CTbjGD4WkhhnG+PstQy0/OT
rQQuTQw0dcMQu2l4gkzWojuKHVlvH21G1+m+t3FL9zdtxq3KvBDPiraLbXUR5gQE7UniiFeR/bVa
hCems1Sd3ahx2qymtwu1afxzfH0Zqpcq3aYB+2duOD4dj3FKY1xuGNXxmc3Soc0SgMmDTF0yu782
5vnEFSgiX8zUR4MDzrAGOenGGVx0Jb50PAwXHYVp/FSqn2E9j2aIdlcb2XGVeNLI/YuDAOpeFeUa
wwnOrl5INcH4JS6jr3VZ/aUQX/WCWnen7sGC/98lPO0mTAlyzRHNMcYwkzLIQIbgL1ud9foxBlzC
IX6A8OWLOprIbd5xZ4IrvzjzYCxwRwGre82WQWi8NHEv1M6BgZARj3eBSQ5plnKkoyNw0hiLReZR
PXO4CBZA/mo8gJl+OjJ8eXFcyncMcNSuKDuhLs9LS6SW1wo+J4WFLKdav+AgWME162oBXfYQspSJ
Ua6rM7s6E9fFdbL6JlpTk+Klkt23VesCAUvNOI5zAW9whEZ2c+q1QKB9fVL3JfvPZmWTKLZ8mbPm
tbbNrR0NBLO1UW/YO9yWJTf7gySfa0vUuUEcdJK09jz28fKq17/vsDXXrJ3DnAO2y9adH/5FJACO
qkkSAlhQRPYuEL86q63OFE8SLSmizUMGEdd2oGVxOf4kxpk+BZc7H9t1bEQOJPTOXvhsGqdNFI5I
oQM695EYSzzDtsVbc8UOXCgBHtth/TGSRuWjfhTc1wR4rdaVfBdT0kWjD/rdtx+9nZUp0CUQlWFK
g2s58t0Wzb0gDICVj5jAAmO93CHfMNc+j55suZp0TDsKQJaYsDaVAppKwAWIFKpLen8fAxBLaloB
/ko/BfGMPqA1377IYPK/qQkXgBajkt4SXtiyLLUJ+L1E+423nNKWQg8zv7jxVhej/gWObUsYOSDh
vvnPVZCA/oQe3TOhmxwcQh4rtDAo8pKfCiAVqDIwJEwCsrGNzHARAt5p/qntBiCTBW0MLqXaEZRS
q6NGHZ1gcWUr5ODdVpKoQLtLMIVbazvTAbAunadlt551XXKsjCyAVBxSEdoA6O/ezvnPHx8nEQl4
vXdHQDm1Km/X9uiIzohoIgJbgQXv25ixlSpn7Y71lyGkqJxP2WDo+jpMojiooVt8dZHqDd8i/L/F
AXR6PPNHjVsDLh/FS5xELDrKvXpigX3ALyGiuqazGN5w8rRaK6x2Zk5S6ugNnX3T0vTZX/sWZnpd
aEIMZAbEexCqdcSKAw5hU/eydynsWS4AXBwsB74hXP0pNvmFNNxfNFITfUTZveg/urx4qKikBXTv
1Hw8Jb3izGEBLZGs0LpbLlr2zEWFZVPcsjrsJ1GoP86+fHORsLFZXuG3YKPKylqpqQlhuQrzetHK
FeCGunUwUYvRknpMFNF0nhktdQdJ08jAdL4f3ejfzZ6dfpUews2juoPgFuj/STF8OdmJDptrUv24
BT4kYL9qvmu39EbwawBe4QmYZGhW7KgtoofvTbnVMS6llhqUR55fNEv8qP4fB18/1wPI0IbntkeZ
LZXJaly50jaacCwbQZg5fyQmWCjJWVZ4buOczqqJyktY2nJlTCOe47HmNpOSyHVSa7HxI7RjFggU
phHzsqxa5kNjEgxRy3WZ4iFDX/AlkvgIVIboZXmRI/zm0lekfkaCUYcC5Bu3KGtB3l38TH6lULwR
DoJcPRBuAvtNYD6BFd6gkI+s0wlEclDuix6gmwceLozUv6WGoITx2qJT178ilIH8rkq0N8bILPF3
57JcxS+zahljDV1aSkMGSZtvgIBIdnbUsF7TAIUp/hi3n4ycXZss7E0wC69AV0Mukb+JZbhxeosk
Xxjz7K77zlu/UBfX9oAhhLpA30670ekG+MUU2X4ZB1+RZTllOFl5GSSzJ1zKbSUavZqQ7Q8CIhBI
P1FQgxONw1I/zoj7K8csiKlu9QTxTF7F1wA+7oC/xDJZis0rIqXv0wAZSOYlIin5oDjdvCXg4Squ
aOqE9jcvL3NsxmTfD8wkLZ8MJEnW8pBoToFgcUtymoCO0wCbRmR7XK66YC1S0H8QZRqLD0+HfZp6
jTxAjCevSr7RJp5dGHiYR7igG62oRg1KsLJzleoSQx7PmfrS/k+yV6IUdTXwjJWsfMc7xxeHSryh
3ZDdSKqrDed4EZJUkhbdjcRP+1rHbgXEmHcDm/jB3aO5xCNfP7TjYnUIhsa7vWjQXa5o2z20pRYt
o3jrx1yWYBiggRBKDzB+wNCfYfRCB30HnO4GKIYeFmqOH/+PUtEiQGKyvYE57bZS8RWOiVu9ptHO
xHPQT9mQWhSnu4c1MNYSwzPuWQzN0VJURuY0n7WcttEHf4mFYqTFS0F+suFWx0KJOTIfM5/spXsx
OesfqDJptuYPa6nmRbGCcFnjFNWzNtLGcmLAiUj0Co2yN60/uFUydtlaTmc9LMvw+HD7JfDd5ARK
vjkCKTcXgo3pNi+JtqdsoM3l5zOEK9xQzNFBGH+GgADx9PzYdqTUllx4ZSmNIJlDh8YF/mpGgtWQ
ghKnMmSFX6mw0ii1F5JcokzUPG7OPJ2PwZvcNxEoe0/XGSeC+n4XvM7yvpQJXixXr8+0zLT4LHy9
8K/CGxER3e8WatC///Upl/tDo4mz8+1iE2SiyhqjC3XHm8x55PvX4evn/p654GmMLEYJ649pN3te
SCmQX8B5yxhEAJGorw7rkyLItRBfYs6DAvK4QHWsVseWKluaFLS3JevMQBKv3mlmg/DtblyLGVRU
TkoXqKJ5J8//NQ4wtOFeNQ1CjnSVXDaXWIFCL6bdQxismLQQbBJpKcejLEvIHiZCoVvR5AQsOHwA
SnlBH0rQDe34vV2B0VE8TkmwqJRpfB8RRF1WZfdHyOHMrpOiADyD+uSBwdChE0UowjpmJeff+dez
udAcGSLIkROtKe+NY4dq++eV3H0+1szaX/qeuZ7jiccmxmOa6e3AgV/Np24C1g4P4Lai9Zdpqee5
BAEu0kCusQ6z6rWBu0xiz3b+vPZxNanop/HBHUMU/kjiI317f0zH/fWGDP2WWjFxDa8hjHEWOmF6
2VC1E7kFsYZXkXdVZ7cc3R2YcT46BwW+IYn+PPEfGcUPVzjrdnEOn4wld6N2EOaUv8HWf9NEtkfr
lmsYDQxNRf66j3M/MCbejdsg6YVKNkCVDvqJwX72AsHWERaOou6Am9zp362LtPoeIQJ55oUOJXNL
tAqaxFE1K4jAApBjcmcaLlupBNasgUrO0jb0uiuTqdv5nuDVYzqV4SspBZFWD58cWLDEJN8jNEsW
C2w5FhdbeziWGPY2N5O4QwqHQrsb4gQjkaWb2p/Oia5eq+MyfDKrK5hoC4vB1RGQM1pMhSZxPgPm
Urq+soYlbsJDd6bYsZln7XpicydVvIFAPqytjAq/zO81kR2j1ZBNOj4aweVxeMEzSmd+D2jbrQP0
o5nxCnXDYqRq4pOVPUp/XtW3eTPrZ5ZBmm3hnEF3T3umAQt97NgJywmpmt6BdsmnbvHz+Rax4Bdz
iuupu883mdC+txqL3EdXh7e570Z2AjHTvoc1X0L9Vgjw2Wh6UDsphegRo3B4O3SP0MabxMjKnhKi
tHZdvLTaxKSc8FK7XTeHD6qDcG3sZRc57FkNUyJ5XFffmtxzvnln/0foeLtLmPqSAqoPCh8KRIvp
IBAO9iPZfmy9Mtlart1PAevH0johex243vuWtnmER89hXAQ8XhOO+HFXZO88ph0bM1Eb+KpBLAYx
b6zOZ8egOCH6w4XIAkuhgcwI/lTeBAyb3FUcIfXzykwfbS7xRLkxsGT8HRLeGqAqWkGC4q1WVyl4
GdnS1J9TSyMSB1ofG1IxAfe8Uck797oglqVPEL/0PFp6yZjNZxnkEtFOVTZL6Va9gPMCH/jdpNzI
JPPORFTwbJg929n1A1A+W6tbxI+hKybD8Vrodofg0daEkkH9ulSqkuhHALff7kOMw+DCVJk/DNjR
UKApmOgSioGIqPfeP+wltudbhZ/RNvGBmjW6hBI2P8v1nkKWNB1/JcgKA6Jl4R6QIBU+Ptd+7MlQ
j3qrO19d+6PsQPRfZlfBs8iGqsG5D9NN3ZR8+uxUoh/bixZDkFYk16LzzA83jHOmnMrCBzUmEbcm
2WxaVQcg30/28gdHT0uD+IgxsygtCZd+B4Ct+gDuHBsiLW+mV19v1LRWXuSjitPeKTDzf1UVZ6gl
GIY4WH1B7CsNUUj3/KlXJBJXbVHdanxbgamxkDuSWjZW34faDZgldt2BzlcGJ9ngoxjOC4vDucOR
1JP/ZYQDFdNzUdZH8VsUeX+eRxFbTprig+7sZlCAG+6aT7ZhkjfGgysxg/6t40k+h+GStbsYPKTk
FMpFqWoAK50cjwKKpMyn+WK/naKJY5s2OpPUwRhTJ96vlbL5ppHrGDDB0FrukRV5+vfMShWBtJ3R
XQjhq1y0Iau9ZLMbW5dchJ67H3qMpVsl7DKABofRA9GvlgTC9yvnNvMtw+vyT09sgM66Bg2kQfuN
GKavfVnZspBmIenj10n0hRmOF/n2tYPoTN2+8d/xL7B/eWzhK5G/qr1X93HfWT4QJZLrDlZXpaaa
oHTuDkzhDsMPtI9/ct1PpDC8ihHm4+dhB3qaIKv30l8Qu2H2zDBETtPrm+NoYTJqTaLw9bwca4o4
7F22QK30dro24P7TBhpthx3cBaxJhSO0u7nW70CPU5MWnwU7B0gCxO9RWPk+092C3muWh/Gk+i+b
3iU22aU1wqnOv7sP42GukcpNwxSIg9lE2I3clY8UwmKHAWkog/QE/h6hBa//UrYExjVwdiW5qWwy
fRHjGA+KRrtdhDa1ycH5NsRNIGu9p1DnjRhVcqzSzfojf25L/o5MVmLuvm7t0SbuqaLe+Tqy0sgC
IrwYXiCpdPsCf/A/xDznbCgrnwDIbayemWhDz8qyJltK/AofJ/etjMXobJl1bS2ktZdlD1A/dN0k
TtzoRnFIOMsRQqm3WSXyTGa7sn5f6dPKuMgFB30k5FL4s08ss5Iu87/p2cHfL+H9g4nIBfUKvp3Y
REOq7G30JWzNIGc0Nd7+nFTtyv4coANcgDIuRZqmzfsVNdyWJIjv6/stn3x5RTRniQAjygC7XamW
Q/fcZ/09UzglpHERhtuU/tNWnKYbZHCfeuc49hv4gvpjJRzRk0lfk/DPjwxp8pD5jN54YX72DkoS
7G0jO0QkCzsHmAD7Lcjx0V5UgeBhXhvny4pqLQTXdnbCGuWwAAAdMyTX64KTDBgPF0VqmtbzGDeW
hOGFhwzYv0sTa3RYpn5bQM4KCDV59JqmKDtqmQiLDjv5YcXCpOO9py2OMxJrpANT/Hp6ZPCa2sqI
O2tiqYpC2vJdgaVnstB6GAcyrOB0KV65F5H96yhkTyADe547aKQWTd69wDeZjldPEm/8pmzP3Mfa
3rQb5V/qytM1+qkTRifvBvU8HXPF8SfU+uvfxm6f9UcWqoZr2CSjFAMeQ1uzaLqwdKRFIljGfsGC
+R6g8ynndOxV5/0zyzPKacEbH7CqFAEC/zkbSVdI4i1H30vklGtcZtzSwZDACycfVETeQHUpWkr5
AALEdJ/WLSghvzlYnYVi0/k6xHUVTEcqrX+pXtQK7+X+HyS/SuQ4J7OzAiXpxcCB8QcCNFmTBzrg
IP6Jl2oFqyVlOfaSW0UPaq+bmibTxAbtvU1hqdsszGTg9IDXCe+g2CWzbcPscNLo3/ktNmvSd9iQ
9Z0WB8zPBKtOhQ2XtWTLlr9FtCFolPfaE5eb71+SiPCrzXOTPnb51kM8dsyCVWg0u1bwaE/DzsVz
VJOLXPSbVWIDWvPDx7lU+QsQfuHUHYjiGk/PIft35/KFATd9bGcMRM4G8OGT/YNF4fzbysSAlhHT
Qz6o8R/8LSqfODaWGEcHuqJJLnfUgGgigbhT+/ePs6g2xdEwYR5kAt1ueHPgpuAP7AukXUqstsi9
k4q7Kf0H8lhQ6nKYiQ6WNknpT+OfzJ+7LMSPLkFyrL2fqP+Y8h1kX7+OS/UomczQDsikB8JM8JXY
ZBbNRhJtwM0D3idNUtL/JRUgiSv2n9W2qf9blYqkDKIOKgfzJYBly6IpLXiMx/ftRvgKxnW79fgU
QHPIVZNRGFyPcKH6OwOWK5XGfGgo1uHF3NAr85O8tOKKVoodL/LTAranz5WmyioWViEEKgGQTQT6
w0wlJ7OYO4915tc+Mj9XESsYnOK5pRnKkadaIBQp5BsC/yMXyUAkCPd2lK6uU7hKy9NZNcB1muzt
13NYWazA9DuSgTwlhupGW5m8+zeEw7LwjQW5m0gtJbVDXJ4VG/SWUF4NTexHPBHEi+CD0ZhdCZtY
gPXy23MFwXh+JSy5JBOfxK1ucd+Lse0upmxksvbeEmcgBY8m8cOaPw501mfZB0ob6gToijnEq+bn
P637BuB79HfILnNuEUIUxYD1obgCWdRNXy0QgHCpf91um+PuBJlGBmsjben4XLCCJiJv1BkgJpfN
rcJP2hCcQOV8JU+ZLlmsD9Pzon0jT/OfKAzMk7pXpbp4yQ+j/fUqLsqT5/IG7RPtRxeEjicyzXuq
oTaNDzWkXVdDLQjwZLZL8pYUvxOao28raRT6JjapJft4lCEewYc46XvrssuMbnMQS6+TOb8udd72
dJo5n3RoF1fMWe4t53rkdZz2luRCAOPalWEwoErgoW7W3rCDvQKoQLcZpjLrBEiHYzsVWcWumCb+
REowQaHIcnlncqpx9c7xFLLxzNcq4q+3bzEBE2C99IuXxocoULQH4nWHJOsqCOSxLxzci6VYODh0
h+Fi1r+4R3Lvq1xA9vA0EH5Avu/U4SxkoGHnS+nBKqHhNQEE6L5amBSpPM0iswRP7LSNMdVykzr5
khUtFAlxJo2g3SbwOBApc115psoX1CiQZRtviLoaOj1EDjuaRmDRsepdpxLJ+4rT+tz8Y1wQ7klh
UgCh1UDp97O6BOWtKxwpXhBL6l4u2yacLpRZ2UmoW8w57PgcyF3OIKdSGbN9L8w4RGxwlkdlkSot
VLnijuttXHJaupgqD9lLxWSdkqbqzabzyva5X4IQzqvmyEq3ryesCL8pjm0sSA9JJoJKTvxAfqVg
8pWBzUKZUTlA97qpxMpRs+kWLRSdAzrF83z2zHCTg7+LYq07If12KsvxkznoSUFJ6Dh3E7iXgMxH
22tuUv9GKhshR/yFEh/guMDupTrbWYVndzgUPna40VXJ/L9E9h//FcS3zykMgqf06y6vV4TlkccS
UeQMHkUjUP0sQU4IXQLm2E0ZQr4J6z814L2seTzTKgzUeRDrzEvW1UD3c2lXxU1XJ46bALvxJnqq
9/KF+Zh/EcOw0uU7yNh/4pA2OlARpXLJPrNritPZkXaZDymxeio2UnDOkrWowAzIwLjZ+pDYFf5D
lqU2Y/983hfoWHO8aXqpw44PosVS1o/azLFP4AeCQI1diODupRvXqS/vBzqUA9BXqUgO5OHN7J/a
eJRcxa/UN2ipS3+aejtmAiW/YJehr3H5nqjj82zNZoSeEUX4zzjg7aNk6Cs4uvXF7kBlg/p8xbvl
pli314YRpi3nAyJta9r4F1klTjZ7XUXUF9DTdGLeWAdV/1nhpPxC7z7prATm7YQazrrZE+7QN5dD
M1P4cIvV/h2lUhUTo3uIdqS7zko5Gh35lYAiRiFiMzuotkLoWOGwci1lTVIHqOhESXVtnT1u7IVZ
s6pjcasBg7AAhFjz59rkKk7NxNyu8aiTMnWOnFpXugtml4OgZallMTbma9NsiypCmP3+g1iNJqVH
e8Vwj57UHL35CgYz9W+astePPSDMdebGXe/ekqf+EoOcWU9fMTkj41zQDkmKzSXIlLsQPCb//Blg
PFhcHD/TT+5Xhs2SJEpy6Ue9Sf+/chc1s/mvWe6C+lF0moXMHj5SXVpCnh29eic64sK8ejTcfm54
ZZeC4NASPVInwIcnIlDslXlZMO+rvGqsXBeHAfk+lhyCcAjeEbKuj6lhllq2qQ6jcFRWCjaRXLEO
zfTL46Ci/TfLGBLVFV3xrrblqPYVHrmHqWTDqyEAKF9lQ5EgJCLO8TKXmYS+Xi5IhNxT+3b6i5c3
PxtAB8pSRPLbKQKuLzz1XxQcuZF0Gq+8bpggSoSlGMcA0+zLnrVYIMDSr2vGvkx1NV2Hg3iO/EVG
JI9FtQQWfA4CuI6Q6A2WDIBEM7b7bgZPkuVMVYsBCPaLknZ+QsbffuUZnHmjP2shQMJ7VQ+0sRjE
54jRT1T8F3h576FGIAkkVVp/Msfca3hROnvZTyOL0uCHJpihyUr00Vtptb6Rqm5os2SuaGq0ae+L
t+smScT3czI/z1AEq1BMdGddO+kwBkUhrZZ//4baXgKzMQjsWneUBMkl8y+goGW6D4FPXJlAO2BP
PY0Fiu5Vi3BTHtEwT1ZKGWN+amydEWD6WEurNdRyCy3XS+0aRdEq9T+qdNn3NQaOIeXZq9qsl/Jx
9K4suQGSPACGGjeAuCkbl52WFmJZ3nCKdeSDsQyhlok15j8uA5j09orR4WFXjk0S2T1MZrQVpvGO
JTszoI3FDXPXYsRxR0/d9st2QnH1tUvYXOQ1E8J2OjgAwzK+mIrxpNa0C1GvkIfTVGeAGcpY/J3v
BJoM3c9/XA6x5F8WCLPt6iyPOzQZIjJ5UzQ29Gk4Vl5zidXuPNmU6EZ0ZyTd+DhlPnH2tLfKCfYP
pAIAXnq7Rylu7qUg/pUyLGK6j1ImXpPnTH4eEZTvRah2G+H1qPQBp+zqC+cvOJyd97HurA0Cz78D
uC5ZKnawhj4389/aDN8H1NmkDCDeuAqwpIJwVXvel/D4N11jWorAgHFf3h+UkKLMaYbExBvX2/9Z
knDYN6mCG3uROyXP6pFbfFeSgPi2PZjong+PgG3zme0q1G/vUjvFJwzuDKFVTKJy2V3qDgY6KuHc
DQvR3a8kCHVax5fR5eqW7gXss9mX3Hc4aNhX6QvNKmWexp0hGRnuKjGWVeqeS0A7ELo0au/FPuZy
L1fFjx6chEVdFukA4WPWRyy94ApksGGMMfsFfFg9tss/FOGbObktEuHf2mFJ5XHsEEAijJAS06l9
isq6nf1YDiGnFulmsbx44XUczqf/8PeRyt+e6mRZvBiwBiFXX2inVUJOu54E4bGx9Z9h5/dVrcvn
BZIKyAxzEWYmC2SWi2Ia8oaYrsnxRyz95DNAeqJEM3dDoWb+ht3reezwmvSRcn4gDccUW4yL9Af0
jzQ9GWHUga5wueS5Xda0n5kn7jxV0sC1Xce2TrB4kVytEphWtEcbqYJs/8MqdrTwNfmhnpwqxz4l
8AExPVmKTGo3qj2CIxLGRtAcFvxTjn5LI0N4l0L0z86QLFmstRA0Oan5Iuz9P8298iWXg/SVdVVF
+qcPC7zhuGyk9qgHP/oYrOg53nHYUb2dpFgjAIzrR8xXrqVuK0pd2ffPWOlm9mqvkn4loE3JKgy8
1vkvHsIlC1opBIsVDjwMMX58VHlYfrvhp65wAWWoUodxPIt1Pn48JKlkBEY7kvs1PQZx1g5TbelH
rHiDRyf+c2AmBpsUH2ftcAvGj8noIJbtY/O+m0PvAFEOWvKjJw0xxejwruYrbMK1bELxnqdkSwA8
Qiz3KhlC6Z2LWhiSMlb65n7Mb2x2i+DKeTpTNIYRIW8JNxhLk4vQd0XxggD2j5hJ2EkPHLj+ZRRc
NiEwt3mTRZHkZP9D2uioI60Q09pJOWce3J6X46U/naoF0XG58mgrnsMaFHTJ+J3OvQDNBHCdjrNQ
k0NlhLumrnMcQm8Dce7z3Sfkfh3EfyY1KjKdQEzGV/kiqgLp5PztfEbJp6IUOdm/Pt+9b5cSCgcf
4LHRLJyAq6CYZj7XvaiWAO2E8T+AW3aPeAKn1lq8QWA+YkxW+W9N0ZAIAQB+9cmIQYshEfLt0e0r
uTcX8XdZyzxZ19+1j0wGSDJx8lI5xZEaLi+X4abh+XbxBtuROZjE64JwLg0d17Y7RFoE1pYLxxvX
Oazh/CB4LT7x59beG0yrB/scXxxLVfK3EAdLQvjKmlFv2c02HoZSg991HJA+LJvkN5Y4vnymNfon
IljHrsbicRnh7QbvCAFsSzKlrXp0pDSyVBsDvvHW79EGBARC23D/2UaOZUkZrFwCLINBepmhorNo
z0XweK51m8oejENrc6hdfSf/E7WIhqhyvC1aah4d1CMILO72jpUEuYISSjbL038rp+R9wQydDJik
NJ9HYn+ktw2/+xmSI8a2CJj1jk/sAAOnHELulip4uoMPUPJ89zzLFavkeSpoHmgHej5a1hdYWpF3
bLb7jltTUFnK+DJBIbxXT+G8OKOfHOI+APuB93hzu8WSFVfeZRJaWWbMGngZsEtUgptklvTN7Npv
hp+0IYMADFj6pLJYzbalE4Qx6D1u8sUKssGKf2BZcvDyvAqdg1QMjUTZFQdVIDnMu84u8G2xG3an
qqa/xLwIkeCWXoEKXMdy5/h/N7jCqczeUYH1AW27Ag7cQxQ092/PhXYJES8Z6wHdIu4lsufRP2nL
t9pN5RD5borXjwpd2/mX3FzJhAQLYRqc2SggP5LWRG5yVgkaxFY0FKO9JnHUIrecI97+Hs45aIaR
vsmL7fvhNDTcy1x/CcEaPu/jD3iFkCLFMTRinFkpOWii3eT+7CMm+WfCspyT+MfY5mhiLhs12AiX
bYrf4PJkcKEK6NZQnQs8g7cduvF/2I8NJhvLWSIi2HhfuLH/I2SycGVA9imeGSIQO+zen2936erf
t/9E/ZIPhQKhOzSoDy6/emw0vL5Q8PPSL0Rey4h56JibtGAcKD/tHTyUDsp9M+Spq6C7LVg3QyUh
MVtQc1j0nRDowWuGmGmsrfn0Y7Jp+lk3NW74gu0jngJkqAMXQ74lzPksE4NieNaajslzBTdKPO+Q
sP35UVLQGxBQ8f3nR+GLorw+D5iMlrPOQHSGJuhMkp+QmwEHuS2tHuQnXppvx7ENmWhlP2on4SMA
8Weyj63JvCir9QuYrKGwZzd3mZtYNFyCPY+Uls0h1dWVHd888gDqUUHWwImWWgfJJHdHOBTTAHxf
FMpYtttFiikuIN3ZyeCD1BwwL/n9Z4cTYF7Ccl0UHeyS/Txex8RAeygquAnH4M2laWpSPiJ7Luws
9qmreceUa4SjXXH5szgFMCudnhAaKuHYhg0BZAd0GseIM+ZqlGxjt1VN+/hB0RAffxzTm8baxc5W
IVP61L+sXpr9CvLjug2CoSPxQr1QuUdf6qZNvHxnQCa9112EDQ/98pHPKMaQXQxBzF4RJr2NP9n9
7uE7abA8lZybucaY1gQBy8P69OiSf+RPdinOBFe35d6aF2L78WlIcUOFFpWuA/E7L3OaNVydBbV2
9OUUShXbVN2gneB9Ui+Y6Vd+KIVliMPth2RWviBl5zwy1luJGp5RYafjkcf9pDffb8GZjHJXXuGV
FOdC7g2XGSskOJxOXzALY2pUMxDNDpbIdNCQZ7nLfl6VzvBO+Vr71VafzfdBaLu1Ii5BLvTPnF1A
l3KMfXsiVvQhLdMq/TqZx0AOCc6tV0S0rLsTavWFQD7b8TRTrki45F1H7YNTmF7dF3A1Uy9gsshj
yksjBlsS0UMr3Ft2r+h3lJ3l+BWPeDbwUuCZfgb/N9kxgaRS1eNXXPYnvLSn+URqslJGsK40YvXT
oTNAtrkKgWHXbB4yVjyani9pB+6dr6GPUYU13gqUThGOJesY73WllJMHaphbBcDdLwMDAduHMxMa
OK/HFg++ZBl1wptlFerKy1i1keLHIWSrn4N/4T0kMB9vvTcSI84F6gK+Qo83XD44KlrgHhhn834S
+cqgwZm/EmY0ZqzPQdqP3HLiMK1jNKuXZAi3Jz6N3W7CGkpk0rE5c96ASF3rr3oFruwwfZ1CgHXG
QfUED8pxxCRB3dTG/rQqD0O9uHAGtlWH66myw4TIiOSpuVlw9b30a2Gkj+FfFGpKIcHaDjja2CHN
udibCpCdzYtRshJx0FS4jTv+Boh2jRuPcK/iJmDPWFL3WtiXIOWSfhiOcyZK0KYXveN5ZBgdMhf4
UJpIvCAliZ+SRg6ZM6YFnIPcpwlkFI28QeTIZOLiUoUfgtlAi3rpa1Bbt4tYZjtLsQFbY9WCvhtx
xenejCCX2Wgp60vYwfXJeKka5RQT8SvjbeXgclDFQKO0ANCn7tom1IZLOWT6RphW6W88ue3qU49Z
gV6GDljYhk+rqxM4a0RklyWo5vLr7Yn2NbCyNOb01u+ACF8enkSD1gLETFtbDYUAwQd2llP83uz/
bPMmIKh9JcyZjSrWYekHkS64AbvmbnM/2oalaIMj6/ySw736+YdwDL4nM1ZE9o4iq5W1RmU+XOQw
y6cB0T4CfKHF4EjnWO7A/wqPQYcCKAsh4uIugX4zdv5dDRipvK4d/zeACnzDUooEpeRzuuEQVeEv
o2JOXguf8f3zyokGqFXJBI438tjQZYZyai4tqa1ejvecUq/DMMpnhWtjFH0ZWD9NiT5Jlg0t3Wpv
db06zAbht3jn0fHvOOsA1E2LZRwUXLHiGEqXOL32wN5GACOjFJz9zWzCdLu5QSPwpVab9/OwSzPe
NIDsbN1VpBrBV/IwdVNfW0G7vXC5epase+21LgX24XuMY9Ki+ICM2dPe0G7ep+cxBFvfCq6akCm8
0aaGBedfCJhskqALx8GaGaK14X4TLiTp+xbBLM4vXBu6SZ2SjzXhVwxdogn5kzPrlljrJI7oM9qY
MAfSArxpwn1VaX8FTZDorIplNbSq+5bvZyQOlzh/hIH+IlPz9sUd/Q9OgtByqiqfn5M3xgw3lgYg
7RjkEppFpmVFlA7Ds3wW4BfXHm06a/4GRRkrgECo3qqlLxCv79J20rA/hWT318Up2I9TDcJ9IO8t
pXBdaZCK+AZkPV2Nc18gWVSGVsL6lu80OHKwoG6W8Xsbtrl03l0nKqAwVOIfc/5/w68CQDun2Fvs
+VLDpAgYTSN+J5ehqC2LJttM22UztKqcu2p5j0D7oQ4xAkTpbaQL/DJXOEoJ7ZA71dNwCXSn+3fJ
H1p1f3SIX3u72ItLmc0gLVAGRqESZ9wGkdQjnbj1pnHumzRUJt3uW9XghuIjtS0J6SiGniuuMqM0
39Reipjujm1pETNErHICPBrNw5Gu7qfEhTYWbtLK0LPR6s6r9thEwDj4S1ZlOutN+FBkmYGpndTM
kxhJfXyEptei8xa7yGsUyV8vcTdelPr0tQ8MKMH5l91B7VAe1sADDQGluTDN/G7BGlByGo9VU7yV
hLsBh0AjxHtIPLdYjVYD3GcE/ulhdEmxgkY9m6b7P6qzdrol0jZWv6bsIrL/Ifl47r7ioY19gxRQ
Krd5Jl0wLK3salvkcvGJE2gf9WrXPyjGv1PnO86jgmcsRA/MO9Pap+8KDRrfiJJ4bZTEGMXu74Oi
p+7/34xwmZLu7hqzUiQhkx4/brG6BbZ4xL0ZzjB38SzGOUA80mOUaQ18NbYq/vRNfonh2Phj1vM1
9S+VOnnzFRsAsM5wXqrgvsRGVh4u4yihGXBCBab+AO3wQasMlE0joaaGBgRZZ96tgN6jyEYF3/xq
VanmDjt4OMmQ4DRdI4kPRWSqqOGVNOlUpP7c4MelCoEazHKuM3VRBQt0B2YaDZwYgF/d4YS6cGyw
RBd2TWKWlRzwWheJJ8OO3S0SiJh8BgFVLiFWymkTQc714Ps9cx9sRuNRPacnGWuU7GWTZzmdf9lC
qmXVnIt4q/UMQ67SFxJN5ZdzNC5xTXsI7EcOwbKQPm8OZT9I2o5Wpp6Mv/SKC8nJDQL07XEGAqfx
dgNFmgmN4BCZfE6lARPvb+lDBLod3pLaR45ji2ADTIn9KJrGu8s+UciHm0d6jBPgTdyYVJa/xfCg
RIABAk55Q/YclvgE9XpQ5B7Bm6bfdrvme6Q0v2rLGMr/wpctsUkw4AAlbeCP31jxypp8FcDwBG3w
YiY4Znpa1ufYZ+gGh/ZmXPSOJnclqt2rLMYnX074hgBlUOzEWXG/L5tOSClhEqNRCBBahHZj86AU
6ceWsWnVQMLbrs0p93h+p7Awe9PjexpPCQQMlqkDlZJSIsbgukUh+drSyo/m6ekz0K/px8kTD0fN
bZUa055mFIF89tdX84zIEwnWmtT+2/fzUGhBTCY/5WFxsKNNwVRiNntwdHi/eXuXO83FnwHYlQn6
98mj7Tw7aDUxiL1bv7Joc8HJPHsZh1JYJbWqt6nxq+GHi5Y5L1HAhJ/c7y02pT9H5LDur3J3kDYk
mAQsVuR91w8Afv1UhVbC38650cYR+Fh/3Fay/GayuNS9hqgKNsnnDpNe2pvK2SdmGB3O2JrTaxTb
8hBafWlCwF0Vhs8QXVfYFE58A0h6kvHECZk+GF0cpGwOsdlovVmCfXyvJvCKKPOrohhWbJiICW0R
1uJphmEHpTMhQ88dVWw/P+nTpwIQCPBZDzmhjWGMwarJq2iHlhCZXIyhseL4HYFPRmt+fYFcanNI
Z8LyzwSsLuPX5kKh7m9JApfUG6HNDmJ/GoPzls73W8qADxjOmW82g5oehDlrLGs2tP/KP/WY9Iub
2+FOVEVgHH/baag9bfetVipkL4ULIxC331pWl8ARKwW6ZEaBv69mjmgbzrpLSRr75iVkpizmg2bj
vy4B09os/ZPPU8qkWzgMQrf817yqF8MEIO0KXcOuglXbHgD1g+QWSNPPHrkiMDo8lnLvOy+siRaS
/y039XBUy41p/qihCKHM333yrCrEYhUbT/wbumIEkPZVQqpeOu4vyriDp9GUISmcNk+loLBIPEZD
0Ryt5wh0sJlSC0RjRulJt5HplFtf4g6xdn/X0h18X9estszXia+JwYGP29pzMecV/W+dVfbqXSvG
KVpN36QrV8NyC2HjUhaqMrBHSn1onJqaDsCDU7nW8xGcV4LRt5K+5JIdIVJDjlVcP7JiJ84mrRTr
DPzxlgIWZePVpQySYf2/7jgBNKFX1Drt0lwDOcHYWv/awbdoO460ay5ZySsJBIm/Kg/9mlzrEyFO
6+akJUtcHJTaOmBaWdw8en74vp2V3wpuqKjCQcyaeIVLSd1xLGHlzGpnYLCdzQ6nQStQRV/frrCG
ysO5iZcnrH8M/GiQ00+UDKkx5bueZAxIDdNb4DnTC+krBkE9x/VDLwDe6z/TswMJJw+pYXowQ23y
GkeOQMiwUr7tgIErWrSVg2Ufwf8MjNIW77h9DVtn3zyrGHWZveAhc7O/GoWuzQEE2Q0Jv6cM2hkE
BC9TIYqONtc501sjHjR8b7erbOhcuUg3UKRBoG2ekP9H2jJSwUDLxYVbI9BBhp+i50qkbq3y7yqw
95cw2x4RaeL8IxYsM9tLWNqi2c+SO1MLzOAhuwcw2aDhGHVf04+ZZlX6CxLzoXOWI02UhlKVhLFV
dC0ZYnyV/LsidM5EmEJX94EKP3hEr2wY/FLu+dyYoFvoxTqOW56EPpCmG6W27A621lsBp54EiJs6
H4N2ctzEKxBsl/Sj6rbX7NQWgwx7K3wCSZiD2BpCpj3sWTJRRmhA5DzBifMvm9yT3pWXgDJy6qZo
bytTVkOv4mJIH5pWV3KlURUZ5rEDFBeouaC3EtVIeohDKI3pFQUk5sTn6E1EERlLS3hYYb2OWCht
mFwrTebwjKMKvvMswZwq4I3MNq5GMaMvMon6EE9+lTWmT7P/K1zu03krFkeGeqdSrHW3WlcKqXKT
cOWmlSgIp+7i3xTU+gEQjeXLJHrZjXH4PukcN6jK4QlYQq+FhSS3oqkYURaf1eAVuujl90S1EWVk
Pxa3yAYY0BMyHqgoBRmLT4pmd4w+za0IXL9FM9mVu55VmfINTNz8LyCv6ZssnynI5A7L1l5SJGBY
qGd8rMG/mHH98vs+utMpKjuDAoHtdQfkTdh+O8ic26uPMdb5Re25pEUfYxWw3E9OppB8HdvjL8sg
IRDF+OvCJrUIvCZor8Olm5z1zsBKGBsi0nkbUkCl5ryKINlSMDYp7qvO0bCdRgMALzq2cjiQNVuS
LS9X7KC9RKVAeVtANYARcY4OVIgoG0UguuvXRer932oxFthMzRAat+TituiAZX4qFdw/o+gXqv11
tiW/aa9i55eQX3so92E+N8yBUZgwH71RyM4nJgSc0JdgdLvA2SxsbuwXt86J6nuB8szhZg+Tr4gG
06bpqfsfhWBfH1E/FKuM3aO7Mem1f5NCDGN+fZ2GeKIIGQWfScsq9X/aTh6yZg6Jyj3B4+5zY4nC
TnTguJ74FeL2Edhq74COqT0GmaSfKKcVlfMoQYjuqF+mxZEOcr9BYW2krKfk8jdvMEIDnZEOuqrQ
wUDHnaq/IbjFii5PLSA34nTTiOBb4vuff/NyAPM8jHWuvh7FUbR23Hkqgqpe5LUBSmnNALIxQt11
P+T6OOM/0wVzzsDVqTD7qVQZ3NtQzWRP3H3VBq9T+TZuF2yvW/+DuK008ltIlbYBIehYVJyz8NRj
DZPcmL64O+YhFNhQ0UYx7PKB+YpvSY91Q73HHy222rNDD+ueiEFUA/UQi0yhsnpmj2H30PsfR0z1
IIk6AR21tIuznYgP8/5CLe7RvrYQO+DzVNakMgu6o4NWA9z1GgnIGe0bXLFzNOGyWN05bAFGDY77
lZ52//hFsqEauXO22bEEq+k4yrr7fYdr96d82nacsCQnh1L6mdROKvmk0jH22eRgy20lzYJ16Bpt
prUK+Jk+YATCy4WEdmMiQjvYAvAD98aI0UgXh8oAcg2VTVkZEQ8EdjYK205agGo+TDNhGD5sNs+D
cpWcyTpDY12jDA2q/cpJiTfiTtsPaipvWlvWeQcXDHIbW4Sj8EOKXMlZoqxdHZZlPXAvgozcOZPV
jmF/45uo++Jd8UsX5aaaWrwPHE5Xf7quN+bBML7cBFTpl7+DyqGN0cZN0shdo2vgUMJUzzMx2zBu
feRFY3YLYuKReiXWPUs7gJzYr1iSfuTn9Nl/QiE/dFkym2NyJhuvlm5CukSry5s6YlNjJDUblp08
lRDhXnd/jiozz5uX1WJfsqGJ2bPRodWWjiUe2v2JFcbCKV6h05XL69K1d4wjCjEGbqGvd+FqgJ9R
A2SocxT/lz+Rynf6XmY2x2xohMHVvsxZUj9aEdL4+L/XtlydRfVVaAy1GU2Rxk66YYIrMb+MHvhc
m7G2/3s4vI0VOjuOnei339NJ9vX99mtaFZ/WDHoE2LlQ1OhW+z8Xvr8y26vPxNLBNNku+LoRpzlz
CiVlxwB/87Xk0h+WjJUwUx8eMmho0HuEYUoEpm2HbAe+B+UnNB+oUPVK3oNtC5wSQTYvK5udbnuI
L0o443Qawv3tVFy9oHS032QXPa/WspwTgBRHtpxoOAmSa9Q4AgpTpgV1iABzuYm/FT5yQCP+yV9P
Yq/LdcQj+9v/ZwChIwvlmIv8HA9n4wuuvE7G+vob6nUfSj0suReIw1u+NkF2kwa2mMsiYm5LtdsG
4Rlz9dMl25pfFYj7fouBshtBOS+hnzUsQOMmP5JK7zMLkIG203EFpOZ4ZRtvGtT5mz8R7FBWmHN4
hbWP8Y17QD8msTDV7pif3y4HrlklItDs+pPmacmcjA40MAAo1rbmwr7BdjBkkZGmnwbZ43QfSKup
+XbXqdRTG6pIUiolOmtkjbbBPt1GfHPHSvZgSNphyPlB0ImQbHyjqxFHr9wJkpUd9HvL3VLJuBZo
D25vGQFGGy9Yerq3cImO9ppmgLMLteczb2BS8co7ySha/I7MVtrRukEmaLBNE5sdj0LOsIElzwcB
CguSgnaBLwfconu213l7nT42A4dh/pKIpItqwxYbafbA83KJNM1OazcW8yEqH4pOliPqMlDMbj83
fFhEi8nE8m4mgo5OUZ9Yo1BwJQ8jBfN545PFXon3Zb9BsLPFzSXD4O4wDq1lI/nd8SB11mOuEy6/
opZp2zSYHOz1Rz8Ccq2yQgyYwxfLrvt+ujTCbruMov013ssDHD4xw7LNnF/XPbpaOqPFVJB+r/0b
P1gxaBIgnke/B4L2M5qnNox/FBhLUVTnpiUnqgarZwBJoYWZtlORdCyjd6eBUeLRi7HZ1cDR+3MK
KEUe0gW865ugVrEvzWa8SKdiQi8T4350NW0zb0kNBqCXCEmEk+i7ZZn7yuVTCQQsPa5LYmN5O/m6
LrAbx+t0OVmqpxa6rJ5Z9EvgKK9l0hHRAurYWqHubbZwpLtERQOhmohxXOfmITgIchdxZZonqpXx
V7BNGKcl9Y8pIuxbi9bPU+u3cyPjODuzGJB8toDLPvKfdtwBo+o4MA/17c1iQdWsZq9repEpfB3/
nEnW12N67D+16nSEOpoh7UaEAnjAaKnR6q8iKpfzpObsRhNfqlHvFGupBZ0RwODKlZSyz3vLkdqf
Le94WPF6M9OvN1+PR6oTk4dAENS2/VVlwNGjUxqq9tSRBC3uIopHWDRfoaUilhw0zU0ZNYHDRL/t
pAkSYgaUB4eJkd7hFNc5S0HuqQJHFTOU5/lHVNKjIPFmlR/EddP9frIjrePJ9dtCAU/P+M9zVQz0
HYJtt2HQGd8YGSusmKmfQvBprt9dxGMJ5I/v5QWrnuGH1QI6Lj8TuacfqdgEmf7/MPuYQjnri64q
QtFfH+U2YqqJUgNiP6VSeLgYAwLzOjj2i/AwKSttZInn7Mnl6s9pAz3YLvrv3OiPVt8IZuzciEcQ
S94b7d3hxU4bqPk2fDD9fKDIUSceYQ+5MGDOank5/vbubVZ5cAqkzYvAzMraSZFRLMbHunCZYFK+
UnqnizC8gQP0bzvu6Vhj6CyaeYSVXxl5ZGfp17ar4urW1GTlSZt8DXMVh/rVazV+N3+HxteFbusq
bnbxJtRHcMMmT8EeNs9Uh4yW2PkDKWDA4lrsL9aFfIuSzFhPXnS+EU/IRlnYBQjZbdn1GazzFcIu
7xtby8OSVAS+6t6TGDMHk06+eBpj8Lmcw9X81oNE8/X9+rQAdB0lqw6XDaXLhOVVw8pOAWHmhYXU
mD3YPLsGp1SE82EHFy1gocV1BQCK23X1Bk6pD1V0X+HYXlZEHaWEqAAAy113LHbSqJERuiGxgtfz
Vr3xo6xsc9E9nxq3+t/QCMcDjEn2OoU6Dmz/DX3ihNAq4GK0nPjVSoT/jk5jb8PVqqp8ToThBlB3
d7WZbvX+n54ZWlUk/I1VR45zOr4kwKeTut4Wj4pAz4w0rshZiygCVQUlIEXVvoRwoT8mv+oaS08b
tVC123ydcwSl0fLcBnb8lC5jpMSJyttU0Yt+ex7dAhpQ1p3SRvTvLxSSBzpZdOKRPBcshIpcpgRA
EOhjbF7lz9YOh/3UAVhLDWBFbO5cNj5RXY33+oj4q8qw+d7siywR+He523YLK/qQo5wI8t0QssPc
fXVYuLurdtZatWcQIl2ohwtxCQCRExukfxBWhm4k/PRR33+n61HqwOw29ukFtvn+ipBFekt8eAYJ
/cTieUnf6dsMysFa4UylQKpHOrueOqzof/wVb4s28AsE6FhoVGR8L1DyD+g/p9O44B5VmlBQsyon
T+lpP7otkJFkVv5czmAkYe0mRRE/Pq5U5bscp/EzVmEiWlJ44yTEaJSmuLr+uLgizkQ2ePbGMndX
OTRn7L0jHLDXU44Ohqazv55g1BD0uWO1JuCyMe+1w8nYf0raso+mDiYZmI0VEZEshKO0er8c/S1g
DblQcljGIXdEjtnOPaKW0ICZnpuNa4BqEc1nNLcFO6KOEPPUBQPhF/LZAYw1ZcgMVfZtQRcgn26R
JFOEce+j0Z1pUxcoIQE1yTsrDdSaYB8gdJeDUDG9yVaGebY9Hb4pOeLFZwIpXwYFmM2+uxlHEpwO
YKda1oDRe+toD1185YGaxuFOqPog7XXOFHhtRQ7JleKfhc6iIBbLoU18gZZpVggiiRXb/96+lbqP
r61/2oLpSY6grJLr1uG70hNTm3UorHjXFVvrrIUkVi23z3VrFo5UeiWB/YX5fJ24r6VcExCoFUUL
UMmXLZaJumXWLbKN72olITPHPwEWqPFQRoBPwgkf/s3/YVu6KWDAzrFv4rwSS544m3oYZ+uvUk7l
zY89X47ULIMKS0YzfD9lY+a/ARI5Bhgm/40+pNf2j9ccJAWCYt8GPQbqOiORPvKi6690aPcvXWxg
/VSkc5E/fUBRmG555fzXRhLczUlRxnU+D6zKP63xK9QVp2Qutsc7nXE++OqXftq5X9u0pKiMgUN2
6eDJsgzioa9d8MnrhkrqjUlidhne11LM16ubqOz8CTTWVLXquGNuCehzoUfqpDSh/R4woZTgtoA2
XZr3uds097/LohHwk13HoJNKD0hxs5HPvpauJESzESkMd3A9yGTtBjt83hu+KFanhpGSnKy0hLHZ
WSuac7elTzlICeVIVwS7AdWa6O9PiJxvV8oBlcz8SDOUT3w6d3vkjTH2wPOK7VPz1wkRfiurczVd
0dbFF3wbDd18yHZ5bDFI4zcmlvtiXAWWjRtOHFuuEYv1apbPMyf6HArC5aTPozr0rBO6fJ/u/ixW
3hLDzpY5kAjw9yclNajtbh+jy1xlBgRc0C8oPCAOXgwBQdfFkx6sCPqqhtHVaeMM5PDzK/oczkXv
+FmPqjuEqRf1sLX+V89JJwpWG9mH5feALxdrYuZ379ayrRUx5nmEOO1MbDeWs9xvGnSWzg+wLDvH
hzeEbBwNpI34NPHGL5LjBLwS2Sjh2VO1nPUVFDoQURsJiWXYksjV9ptYfy0HfDwTqhiDevLw7wZj
GjZamkOdhCGN+mjQNYpH56lhEXUsc2aKzZCXQGznwKIMNU9AxhlVkd+JTV9psuNcvv8qwHhAnrgi
aNGvGxUgiftQveggDp5zZe5akUvTlTTvloRA82lv9291DXjEtEaCE0qs1Ln6IURi6PrTmnUFtRjT
K6YwX6bDRq1oTz1ALPFQx08lYpza2ZUhG4HHGSDPL6fOb8bR5guX/wFpToQcRof/dRLjlUlPvVff
F80CqKdKmE2UH5IJKeYet2SzuXf1OsgH2Gh8LKAX2H3rAhYnNER0GNdnqiz/C55DR5lL50jyaddd
HmPFq/71dODdLHDxrB5GHIdJpCC5iqPQCprgfHA5NuhKSTlgwLHxhkMCZMCOTEwaj6M/rfzzK+O6
w76unQ0E+5uSET+5pik+b+cbkBHASz3oU3GQ5zsS7pGpc7wcVedFBnSwdBbr6Lcl/+Jx1Cqafr2e
Ylib1OfDYhjrWdS688FXsVgxY62tEGl+muaZe6WeVbQAHvFPK45MlpJd93E/9LtWzI+E1zEFWjAX
5/my/xzMvt97Hbre69+8Q5wXl9JZfNGhtLR81zD3cfjDyOVo3LR59G2GwsTPEuBAMUQbDwiZ/KG9
6lBllyr2wEkxRvihBjCwNnaZtytDZ1rQaV3wMfRSiOmiYiG7gKcbEuCFHg0skibGFOpAWlqi4bzp
EXhiMfmMzVJ0ZYe4ySzWb708ufH8FoL3klioQHC3cI0W57efV57ZSAB2FPlgE0/HoP5TAIUlYWuW
g3hWqJuElRURbUpL8PvJvrvvtqLIe/MRLjq6rXf9pA5qb5I2llDKKtKTk4UjPBDPAw01niRsy3gn
7r3ONNO6VWeZANbBF8z7vTZk7wznfLLAFGI2yW6XL1dhZ8bEttxhL72iP0EyFzjT9PTWcHerFNIn
tLON69XipfRoXB4m8tUpmKPqW1lG93v/mmx60NpOUAOeY3+c5IjwUMpH4bAr/M1n19X1J/uJvl9z
hUarYEeUczfOBxL4ExJVIoSPTKF5as1W/zwScexK3b1ZqBQIIHUGJI9lG3I3zqzpVtTiAXNOF+IE
J+xFaNIycuZoYHnxAs+hXT+O+l/bl0bZyhHf8xjiEcJHG4mRxRgxjrcp1gnnWQiGPl1MUfmihbyA
fQsZ0DRCrJXdqlaD1gi91PE0ZCVoB3tnlNN7/XYloa8ttlDuHpibuVK7ci8XGBNRES0gBPDqIUJo
TnQ1790GMjBK7J+EqS533fGhw1U3f/FmdHmPvCIze5abJoWY+2Lr2LitQli5ugCPH/iPcE+cPdAh
cssmtpLN8PUR3yAMsq0/2G0FPv7IxKcapNVg6AaVc4yAiReV9JtBvcdfX/BLQIZYIGVja+iu7ktq
aedWte2gIsWRqPduppntaCilemwES7WHTlc3sqBsDfn3Dwx5LfNrfma9T30lkC6VeTuPWHm1mvJL
BKOhGZlnUAT+avxNf0P6cx63s3LMmGM65Zrhaz8RejLA15mKZcztJPAGYCrYlJI3QfAhw1EP8yf3
Kcp0KxkN9UyV38BaoSmUWpp9u76TQkREukiNbqDEDSOwkBx+BxxyDneDH+Gs7WG8Q7l8jvztp8Su
cYnlWwpsb+9q4d6da8CAsihtJkbr3EFAodYbMFBGyUKUSD6+FX+5OWCtRbTDkk+GTd3ybdJOhKhl
odA5221Yf6YK2WkpokFCLGJX0l2joXuHmyPzaPdCF/6MR9uj0GjTAtCMVQ2pCC0ljsVILSxJRlbn
BV3lcl6HjF9izWDLcg0WjtUwaj0TSBAXBErY4z+7ukA49ueWjZbx2v/tQraANL9M9Orbn39bBFow
hAUhSFmixIkfXRJfSBOYZ2QZ0YuU0QMnQU71dhPRWBry2s8xAtWWw1KaPCJXOJHGpKqtkizaJ5M6
1FgLkHjH6XdYXtgxpqhe+bNhgH93vk40Hd1ZS5HnD9tdkBqQHliZ19/2NBAZxv7ZqRmg2f98ijh+
d/CzSgPsH4NE3yUKWxmcEUdwT86+lb8H84yAgSeKJDEC0qzJTylmgktkmIHCxvUDNZIoVLRUhcIf
bALfx8osxpgWlHigXdYrmaNG8P5SR0PjVE7dbwYLJ6+vHGxFjpEb/3jHsimhvQrF7ZpfJ97BqLAg
KX8CWiEVqSU3J9LWLKA1I2pB0kfScXrEzepFw6jL1Dm13ATTuF1tnWQUfhWWx53nTQUgEYMY4nxb
eTtxSFOAMuDbNgcU90vStgZpdC+YgCkjuJs7sllleuDXS8BrSDEykoqcglGxE3kjzC7kKbzsQRak
lFvGPAl/oGLpmQpBSXom6S6IeSz2F/thHJO0O+Gwv+K2Yg2BATYqscwKSqw1+7b8TTj4KNxh0uHD
fPki81B2gYbe6/rroJ/rpFA6FnKsLXBSE1YaZaELigeuGp4f1crKZncGqWf+oEMBxzkEeymnfy5l
f8ZLB4bfoIAN/I2xrE3x9q5y5FK/pKiUHfokIsIe0x5VC4+uu5T/JLdXnJ+fsCPI4v5gKZb6ovdn
NPnlbojYTHeUaRlkJy2jCipZPb29aRU1acKrLuURymuRwXh/CyoPtdUIqAEuZRCDZlWcM6h1hfDd
iCmzuXEu0BaD7AhKHc2UpLtYF7YxlR6F2NyqhnaykbHJN/PzEGht9neap+v22ksyrRmNFOCjZSjz
eRYxJaNkDWi5z/ISuRD6Es/aWk2XJwnLnB1eI0Hnzyf6jDllys1Tt+9AXomlJR82TML7fii958CG
qbI9tavoHcOBUSHn13IshCyF/Kr6rGGm/j5uNplGhPIiF1ftq8rNFRzLetJnkkfkvYZH8Ps02R/6
TEhi97EvMGr6KlhMIBmb+XQwaCNIPHwWPlNk9rR78iMW8kQZ0R8yfe41twlsR3drgF0kUB0Xn9c7
gJyItdwD4GXcicXjnaeeQsFmqErLLEaTdTwJN4JeuMzJRdfj3mxlD09qAKuuqXnQLS5UqAKxnIZ3
XVJWcV6s5R2MMn4ggds+JApzJYF8Pz18XKWq+X5vPbLqGBFgmdFaRzpBWaTYq0pGijcAX/40FBUh
Hp4hm8e6GwcxzsVOn5LeWNuMbBA/joDQh58RF/9FhhPrgImn6SPCfw/EtLJnGOZlIr/yO1Q8MlRh
EopuG/q7oIWIcpTjgpBvmMEHV3im5TXz6i4ZMvu+/vQMBMm6WofHrjzHgzQdhX8eZlZ5Q8y1UTyQ
ngDB3W0M+TqVaG/m1NvAVRiQesonLh+vIIzjcFC3dbLJzuH5pw4EfKtoReIz+nmqoLNy/A3TBpnx
1pX6TlLqD8j1pfngkZoAKSTcGnMYk4t4YX51LYX3iVUGesfVX6tjP8ooTzuDD2oqho/fPnODLVfm
F61onPtjABQOTgV7A2xXReQbESL1JTwWxOY04vtHooubpUqMVxhj5Qom48U37w3ITCghjSALoTxn
PNUoZaLCzH/J3cJnidoL0yrQDf600FKKxDqENuPL6UbNgt/u0wqry5hhKsgp+XtBdgfxfufr5dZV
qVDQwb+HPluiQjpbE8XzIU1fCNyHzfPHYM7559UuHzyGpkJEGwT+m9fpoF8OvIfq21Zf5jZh3AR3
9il6g3o/upOjVVEWTQMTcK58WBSLOSIlL7eSzqJZqmPeSOjmOmhjktuvEKgNNGfYkb8GxhZx+gWs
wRZIfJIMc+6SWFPt/bhFrQCyYtQk7QcutE4jWonRQn/FDCdbfeUXwCLJm0OCaC7yTVEd01doc7ZA
Sh3qrZ9xhn7PJfKUHsxV1Arm4DKfgMCTJktJuOlV4Oyvn+u0IwbRT8wrgBCKllhziOKUIJ6JMub5
QsDEMc5HaHNzuxo7yC1/mnF8MGWBHZfJipeFOaunDGbqIpq3a5sRwEdMbXf4/AcKRAHdJL/zTjtL
OFOvtkK2XfXnkvymlzI51ZYeVdyyIShEuugwrBNCNLqeJLBaoWpCNe6Mxdt5REATMfHETMWLVBST
aLq043j+TAk97CvP6DdK7KPH3HOtkw3Hj26Kdy0q0Wqo7pA9mFfFO6qcss3pDPqGPjTccvoA+9q0
KrsXU1oSsi1uI8Ro/zQ6PyQojehfTx4sHEJTng/eAzZTM8vv7HsVTgay+KjeYcwge4QsKPUYcxbU
iFisL/gbN7IM9ij7NtjsZuIPyp324uWV7xKgYaJiF5Ud1sJIa8yD2yAYDvZQEzxKtwq9aIzJF1h/
lKF6uuvARJUSdU/3kryiyj+CXXRR18onBQj0+HPOTJtGI+8oB8Py0VXleADQ1wrnGcrSRd1Rtkin
xjbTnN9V91rvGHAfUogVDlkP/MdkOtNfzaJP7CaREWxqqI1wVrB065sApLe2VX5GNkcqeAdJAF0T
lZ9fA7ioQcLf3zaqiD3HJ24j2QCpo5hsC9fjpBu2SJDboTPdYli0aBU1NKfj+knxbJL72XRd0pbl
+zQ3sThNSjz4fSuwQp+R3yOQYGzWKXSuOWHJsgs9ZYHbPQuf11jN+R9EunLAZnbHGbaRgHabrx8O
Wu+OFND4LdgJgJ8FGarlFTV1xPxTwoLR1V670UpRQXlThAgatz7h+EgVCvxLpJImwRsLHvHwiKHR
MmiZvEP2WWB/HDNBSP0DSaUJA5LDmT1YA5ehOcCoH4tbLJk+hgEUlTQ3y7CVolqDBDdXE/3iIw5m
XpJGDBhQv2ACCYO7tDEaU7Fl7rl0lb1g5LBdYy3jLESAW+CnfZNfRrnXHJnzoZn+91GHYJXcxUKd
pD+ysm651EJ15GCCKtnXCG9wkWqaR3SaFKdHc7ND5UPHmmUdX6DgNy/wisCa6pke8FoD6OYF1jbP
/xG50RDHHzwWii5Lj74gLsUyWEtcaQpVm2GEQPpxBl1xbZvJPF2zb6/PW0FTld8Ns72758fgs7rX
Lb9TzrGlgW+wjRODZA+ZoShVtwCY51DY+N8zLDeMMl//8jTKonKgNQsfa9ZVr8qvwKeV9746hFvW
XmRvSMsKXjX+qQL4RYGa+tpjMyXweoEzg8jkZMsyNAK2/EKUFr7F3P0wcXIG0ZwG5p6UN/NVJi3k
ggzkdR7KFspjbEa46+nMvrkR0nYBrDydjJsWuDw0MVOAqEbhQ34GLyFRBgn9ALROoxdldOr81GA7
XLcdS5b3uKo5Zf95+pLntlJljiD8Hi/eQTPIV2BH4fLxHNFu4iBh/zhO9KEu5BfphHg4rVS+zBhR
2j2YFgP3wOPxhNy81jog4VOuPKQ8Wh9onCiptnMP2e7/CIYUc6GF0qERIEkeQjQNoq2Gc3wjQ+CO
oe+hw5W4oAmQsXT+87hOaxIbad9P1Vurm7jkaQNWJ523NQ5Kob50G3cfLrirFINijTSEMghFWFKQ
rwaImf6VQrEgRhFSHKt6q80VeS5kR+hw2e+t1ArVIzU0wTsX4dNvlkxxQghFYB4Wn+aQAMZWYuRZ
7EwUmhYWCkvlra7I4hgz5SFcjWiY288A2N3Ma5Vw3cIDVpwrx86W6h3RlAljwIW5emHKW2FJegbl
lifT0iHG1Fd/Xaw77KqEmfDjp3Gova2t7XU3L3fAOet981N/fyMzgRBk80lwqOpOx677qZkOsMg7
NYBr8b5RCNB75i+4nR15ou7F2cTqFJIdJ30iaiSSHj1zE4/ENpIDrEUaVeimWX+Ij57+1lb0fS/o
4eREZVpFS2MjO/7165QUzO/PJuk1Bou5W89CiHBj1ooeM04yrl9Z9lYO/F1I2tk1OqdW5Xw9IX0c
qHKXGQg1s0ORGGfCsf8FDliuVQN7sIkXBsQ2iWzqjwVYvaHfAlduu22jAtO5lK2B2w3MAuZ1Ra3n
Oadc18Cl0RUvHez5RBzDb65RHN0zO20xJd/bcmA4Qcch7K6N+UDuV1pHuhfLLqHQTwLzT184RVR2
uPCOpXx3g54jgCJXiaYf9LDdIHT8Gdcyfuwlqj5ACc+XZWb9qyXe9sdKsfcECwrq/vs9jIybhzLw
yw9d/jj7rElcdmKXc3bIoLmZc2jQ106tU3luAL3qEKzIK2Trj5pbdXXuKFNRZKfwENXk+OGLpmAa
ub8CPkc2NIK19hi+2UmyEfg7/TfT4S1IJZqLoly2frEqBX1xRzFfuIapHKzaZamHGIE9jWgQ6eMa
aIxgIA9JqcqDxsHrShmta+UV/gAQJu0ZHnbBpRX98HY0esQxiYlouMTPzZRG1S5ZYzG4d/VtV/B/
YezFfqoXFdeiYleOEFPr1GhOdh89Ly2KdMNvaCktutCI490mjvuhayoW1sxQrEAzKgzfH2FmYHbU
htuNGUoxpSRQvsY8TMSo+nSefSVApUnE2gFynxE0rvkxdNjrRAloR9PMRJNhAW+PwHyHhBsl8kTp
yNeO9/7LybjE7nyQucE6/4vyoioFg1JX+LDrUEayN7EGM8JaNRMBdjhR/yz5oc94ky62UCSXq1az
/4mmmnXV3/emmU+YOLWA2hlMEcQzixE3SF+LpMZbzHOg4pb5E5c/BnSVB+3ewWGUjR/pQVfpQuv1
p27N/TWwg3J7bub39DZU2ZELUNQYsm4T/OORpYXc4zGLTfbElD9SaAEAbYaqasvMIrkeZBeuSxFr
wBJanX1vAY7jQU2fmYHR19ncPC/xNS48pTKWYQCvPCvKw1UZ/LZba2/WoC20YZI6SY3zRBUzACB8
0kl5SHNNTID80JlsH/XFZzXPFZbTy3sfsOLWC/ZyxeCc05XYaw4HMcGzRyzoxLhjXb6vh9229d4O
8vTJY4RGTHIy0p59kRvrq4QtHTcWhPzPWwIp5ZiuUz3wwiGRJz3ytf5abmm6lMXDOQFG7mip7fTA
QZtldI7Zg7b9new3mpdFMYWzzVbXPwH9JcONqBko8WfMTgBWJEt6N6bvZcJ8Izf0YK9YFrf+L7Uo
W8zB/a37dIcyz+mD9vKq4qRm2RZeXTXyc4NFh36T1b894ZF9lQC59/frdKWGmTwi0eSS/GIBQd/i
CNDDmMMln8b6DcHpoKlAtD20XFr3Tv78zydq83QW4an0/W/XggCVN8Y+OrYZZiaml41haWaBzYVe
XtkD1VaTApzx64ul+VutQenQ+fQcIDf7jRbdar9OgIYy5cKe/brp2qK55pG/OSi5snM9Zv7NUAld
gF3E8pdvL4IUjBrb5yVtGfnboKfdLQ/N9prjFTlTI87+7MI6PZq/rXfpOhpV+tJDeN/OaQsFAHwZ
BEcLRLaTfTrM2L8j7aeQX88ZBtsyiKOkg+FD58U8GejGs4qGF2+vifQLuJeRNBO4mtCIEOQIenKO
C33tSpE2a91DFpj2mUxmbREWAbaQdRg2K9X73n2kB0dvmX2C1BsY4J4Cb4S6Sh3SUfSj5X9C/Qiq
ukRy09FU9D5NI8OIlgNgGTZ2MnKDYAfutdRJObHxOTgEPPnKsZJhpNFhu5qtEGsgMgS+QMVsJBeP
Bovm/6ksiXKaRxHhg5ViWG4f12VfZFfR1cKcjbyIbbSDoDiV9q+XDxQG+I2m+Smlx/OWPdWMr1nU
9kmYCgvBDqywAEvtMzs+zTQrU4k9Jmm+p5b9I8Fdfc84RPPqhRfJHgjg7dvikUD2K9FG7zZ3Yq4T
CSDrMumZxaOCCi+izu0PuG12G5QaXx4r2R+czAbjfwbxeWtOfLsZKBtwiCMVm1j/8VpQih2nhR0M
Q/RGO5EH96BajIRwGTY7jZ0c7K6qeeh7pRTSkBOl86xDbcnikeyEkhHDrblPrp4L5L0ItsounE7p
iGrfoMpKXrEyvd3+U23SaxUANgfkQoRCN6LB9gfRc+1GC3FOFy8Nbhjz5xJWr4WxU64ZtG2XqWzX
Z1xk3C8pPlONSUEKPiGxoPUVadZbd5PBWZKbifFe3XHz6tHMQ5LfWC+eafQjnigyMntl62aiGnoA
/GQgTnTzvUfm6mlfTOvXngHHAZTMVzWN2KiIrT1pNCZiNDRXRa4CG7GcMQ02OBqYti1z57GllAEi
OO5sZ9E+mW6c33XhzrzNwDAITpvdn17ZHEvMuf5J5DGyUPjeL3h9s0dzgFPZCz1P7ur4DhYgYO0e
5ndDq0b4ZhPHapaG9WqqrKX6iSYoCC4xewZeJRLz7CaxZimdQ5g8svp2JoVlqV4k9qNoIbGl89IS
ZJiAaB8meMTC6cgEWWb75eEv3QbnVfO+TEjUG0MfRCP3ONKwsrOGj0kj3j74o4Y5QlKm+BgNFvge
nfwTXypwE4U7pQinG1PU0xER47o9fkWJsA1p53PMlywGNQs+kKFMimeqAl3bAhDrLLzhVvMsGPM8
DWTYkk3/0VCQribsloxKkmGqwFyRmRObPLrsgL5VSHZridfBOcZNwr9bQSVQzOqisdlIZCnRd1bx
gFKfPP0NhraovtPImFJvjoo4J5MxlJhm5S73aAUQQRTY4/hcZRx9S8wiJ0fISLc3862n7hS8Yq8C
LbkjB6IBFr/8oz3q21c+Lyfs1h47qUpVVQrIxOVaxzHHgkZgV0nuCUmxqSn+10vuv3/KLiLGAg9v
TpSmKNDIh6o+AkJr0kvMT5s3uRN4nUUxK4xvybqN1D6OhsH94W6OKBPBSJfy/k7hA7rVr+rrJC3T
0d5LJwrKEoWtpLuKiRDeEiQHqRBe8QpdGr3m1YyJcXZ5Z1x5C8ZLCmRqdlTv8ixy24K4UxcJeNQ0
teD1oIyCr94hVJ8xD+CSJXKy1FuGffZOmDFdZLAUe6w9xFAIZJAfC4F5GBvfLwq9JYB3aVfNsu8V
rXhYMnJHSTfjnvanras0XakghU7Qy4Zdp/anaZiB625xI3tFg9VeLJsTznx2lm58XGOMsx+9X0q7
48FoPs6ISO2SCWiDjnndqZKsZfm3BK7DHza3j0JgDozyEi0hwSVx50tTbxWQtL0/Z4nz2Uu9FDcm
gcDFskPdvM5mhg7OFg9oOf2xKvFvaiAXXu409ufOJYmNI8ojr7FZcQGLa7bl8EgzDB9SU4hahdOa
jHFfJ2OPd1BIjM2T8WkTR5qy1hovhOGwMc+haSs1CNFfWW+eXsWmV3ydM0b/ja15YaBIFLYXXSLp
I4NPtfoRlmQ2VAvwA7ORZakN28rYfLpXc3jgEmI68F5DdU7yMrgVgCj7/CzbKAJ1dBoX0WSdhTIL
O8623BwaLrOYl0RVKtlboY6O64KecnkvDHSgENvjdUNNQQZHlPMTOugKORwt8ZHCvPKJXeVbwpA6
528TkFQJ+oOz1TbFsxBgW1matBKUW8fe4fjxVdDMoTIKuZkPJHUTFt8MW7DON9rm/Sdp6lfkh70y
k5xZNGrFBguDIKQr39T9uZ+/oSsSJaee53aLc9WZ1fE29hurR35+hXBChFRHYIQnqX/Kc9sa1lsa
SHJ0Clhi/+H3aSj/RhbTTg3MF+PGERa6pOXoz2ghnPVfzro8JvtMagDY50aGw26TrH8MANGj/LRG
L2ELc2XSxnRpB2RTjAptdQaC3b4L9SuzPTbY7x7+BSqlN6b8ZGNxfiIGMetpFgdDbaexLst/k5Uk
TU5kQEz9KGYC3CFCmCnHCgHuVetRK6sOaoYjl5F/UXJXaIVHrvMkJjPBjkzGgtMPg88+M24ta1qr
dYA1B4LAzbySAtQfVmRlYDZ0bc59MbxOPG7PpPvrKEJXJEMV5OwbrLRRRt9z6ueWGWgQSDRDtf3o
SUt6meacBa+AZ4mRC2DXEA6dTXy+hlrqqsWBB5fQHaZobWEB2NEssJbDYjNBjokODtDCHu5BCCcj
zUWb0+7lnNx92agTTSyEcBfuao5fLKJYbjqCEEzfc1BK40k3/kDx84iF8aHTvWvaKApphRPqNMYk
F79b8/tLa17PkWvNv+iupNFKByPsKxyWewGFS2hSOIrY8okSjpcREidOmvoh8xZHx9wgx4Ri6qFT
ewNY4xwLYea2k2not3weuDUZRZRirhz0VwlRGhlk3++kzwNskTvpW7tKvOYDkv7fwvPaoOUeDwp0
aVzoj+vT6z1jNiitHaGJZD/A3Of4AoyDJLLmxx2geTIydM/7P0+wCz7GdPMuBq/mPvxKzQS52zeu
CeBtFV0NL2Wcv7kVU6NKKUBWixMI4jXRDVOkA1RBSTR12HnP6lr+dYHNmh6nyt9gRB1HR8ViXa7E
riS4UvLQnlrFPscX3StvuN1ennJ0lXAuFlDp95zXedXyod7cxiD7hiomNtqA22eL1RahGhiLxUzq
oTi8BcWBLuil35Wn12GBZBRlfb81hCaINQ/rERlxsu4jho/lCJCGtjzQLId2RTX+GHT5fihB3dQj
ELt1KhAKMQ1Z4kSrWAnoXIdzGxtWoU79K34JBRHsCfgZ/nXKLqqSAcrESX+HsCPNbeKmmVIEeAKw
9HMoBkKcwBrf2g82kw2k5vviHY2fayWPYQv5Jr6OvBnTTwSXiqLiuC3HV8b6wFTCJa1IhuT7R8mm
h0ELWYkg7SmhhAiLgtDqsAVmqywOJcmybhxaa7XIuZHdc2gQMWN4eOcaKvAjhIasr82zJY8qd8fO
Ub7PaLC0WxKdlozji2AsIWI/SA1peA8xfZ5Zuu1sdimInm7LvFm++qjxVomW8u/JiX3cR5+pMHc6
lI67QqP8wnZ54w+2Urj5/BgHhZMICaoXz295Or3b9sXVO4owt79k1QZrv3D7wIgmSF/2iN+TiPeT
VKSzh4oZyWvkNrS2r5tjFGA2Alzd7kwBxU3olBB8Mmc+HAaThrtgE5e9PvTVkappyvlNsRh1AOPn
MIwe1shBAM+dmAs0YYv2iYju+0Vzygglf6QVQZYqXYZIleexLYKs0iSwLz9aM9P5+xuMYIIEvgjX
Q3L91G1p+TvzDJrHKh7hC2CJbp1IZTx0DkdfyY9ZCz7Hr2YFRv7f4HrGw8VTQxG0j7wOKF79Y4nk
8l40NcPruz3B1G3vOz4O4RuRe9+t0EPkZSHQGMQMMMV9OhMj84tuSZ+WD/BCWaCSgIc6W33WTFHg
FUXyMb8iqqxsHawMF/sKAOZQYqURERIqFgqfXoKqkkprxWRsqrhmvvnov27r/5k5sPqtSPK1nXrJ
QVO4eruOR90fQnGDXwjmBWh02BUW3KIduvp0n66J8cbuG6J5T7q1IakKhHdUONojreo0HPGQKm8Q
TlIHiZzzRgWFfGVAQotUvU6GpB1Li4ysYdRnwhfi6iarAEWhiOvUwqOwWKHGWXC4Gp2EC9aZa9HY
AGbTRj0FU4jsw6SP9aQareFMuaXqSiN7g/D6RqHUX+VPdiZ4TYCPg7dgWhaIb+ev0h/EIB/NwpFx
j/BfDlMjnogJYxK4kggYBLIw2V9ajLG+qpnWVc2uuYpeUnslI97lDkWA1tWPbAym8tx5pwHjN7OR
18nxtkPrSizQBQ8Ts2bCzClRuPd0oIVpFg8ATIGuF1JgGBkkIVk1U/5FPK+8s5rJPf2Qr9A5tZNh
d5pB4e5cO6ObKx5MhsPNGhG8MldHNAE7Qrn7LpHyHdpflyIEe5o1pU5NYVYaDGWZV+4ZFHYhjwWA
Kiztjslp0m4Yjnmh1B00EnDxF5Bd7m4Sbbg4Z9V+3HMr8J9M3qwGt+BWfBS4taZbqdlAg37ma/RQ
cJcFQwR8LV0NBMByzN2WMyF0hDHYl/06TrbXnVhMRD7bsAp8DuUadsQeQ6Ax+jNlgS+/0G+4CKmn
VFZ6M7UmF5s27WHScdZ3c7daIPUWyNvo0Pki9oeN2c2UFkQI24TG9XH+7NyCL/20R2dCmrigHvZX
r4E3IZGWKGpe6ApqinQ+TbU7+AgMMNf1jNx3GibOinU9VQEEUPRhZD6rjoFjH8OMLv0wEqvEF7Q0
S+o+gusi8Jug+QyJ+l0Tztl7B2HcosCg/bX/URnE4VUrOrBilQVFeiq+NaOvZaUoNpeIAn4FwsTs
yOdfux5PRF2KWfKYrwzlpIKJwFiH/KGY7dzoc8IIyT82L1qJl3B5UVe1Hjk/reVUFtgzyJP8uoUd
SjgThJSt10s52+i/6033eWE66m1ajsFcw+5HyNHcJ4lnjHjquaevxxfJFrW7MSAWQ7S7pVu4oBEe
NV+V1m2c7SL4fMschc13CF5sFzf7MV9xR0z7fK8DKnfmSfDZ+gxibvKBAAq1L+PgxwIoQyMZemZS
TnkAnWQnBgTV/AikJMmW36sLpHs7P4fbaWEGlqJEHJqSbpzNiiapULccqzY3UE5zgmqLZi0jwwlF
pKmjbINeWRoqD2cBPgsA3Bgy7Nth3lOmvzoWoZygSQOl/Pd3TpFl8/CSb6/hlqEyHqsLbz6scEDr
69fsA2vzNY5xV+XRDnzoLQLRMwO/jTJKbpoq0/nXR/LVYn9eZnaNipTMnZbAP4bVA/5TJ4h3hjrQ
cUGfkdikc91v56Qqgp8d8rcrF+NQoD5yQTyqObs+iqQaWghc6npb0X2Fx+q6Htx/WhORemfpQpL8
vrxXyaEqTZYhO42e8mmRRxp1erhc5aaZyYbPRupCtvkIeWcFJiCphUsvAQWd+JnS+sptpVDmW1E1
luyXEwKJDVTrBmQRFbplZrDxfeQJzzENyD8I9pOm9feqP9KhQV9pPi3RGesu+xAP0w0jEAuZNeCp
02b53YP6aOCK9Sd7Gd5MJwiTPwnVqNwDhUzHOOFqkg/BhzSpokuDDTmponeEtimv+h1Nk+peBY9m
/darHUrpviWY/yTN2jWhpP7SIx6RLTdU7py+fHlx0Sqv97ZpY05ZYAMFPAWVItirE7HIAUTlhRRs
RLr2V09f/XMyhq0PPGNMsHWTyUklOmHiD0PQIqsdzPQRwlL0XclOgf7yh435IJQeFZ1eImzJ/ugz
87w0qq8Ah3kUyoYcKeYHx1n/Q9vWu091PVbHShCY/gIJDNUS2QfWSFdsv/OyVdsWQdZ+soHEPSYF
EuiGsWDGsFouetP0uJqQYPbpTqdXpAWaTOQ+uGyTZqzOcaRff5jtJ8TFOM9EGs3yUNHaNlezHz1Z
Zjqv1JZGxp5pVyhgZF/994MsKFmjdLPyey1+a/em99yGytcSsB/Z/eX58dUVAVH2zeuW/9g2DgHo
R5AofmaLU0IVBul7LN6BDiaP8z0s+8UR7/R/enzT/V6JHAv2VUEFF/gSoztrPw0fvgqAoMZH0ro9
GzIvesdrD8FSi4uu5axycnW+llT4/M6kmg5K/LTksKb3IDTyenbP+iunSrZ2zfFbha4Puno4q8J/
t+9MBRCUGrNi6FfLkAudVHXp3cHCiO8vH6POY9gtmXRO+l+CHfRyl2+eKSYVNKkmypUiyb/VeY/O
jRmnfWq2E+FefR5jfEkZdHahuR0wxjXv61aKZBXb5PsqO8zZ2rdwowpBskBEBnfys2pDTfH4AuAx
NBIJqm+f9ZgFdvb98GiyivITrenZ84XFAKitEmJ70vivstvBF1G/zeg3F2wrZVzI1T6gW/TnIDT4
dn2Hlp0QxBs8hZg+LJTYRyCewCuZ+AOiZGZLeno4cu4I1I/LGC0+hqffv5oO6d9gFR9Cmn469MGP
WSh72jpbXVPGcEz+T83LqOVTbjHt7ctVQkE8MSyprGOpPru0dmoowNLOh447W3cm8Q3oRY8xoTc+
dJ0xHsSwTPmLmF1QBH/eZUUVSCyWgmNzp/lt0ui6F2vXiOF+UWLucbj8gwH/pS0Cch9EVKcK8lEp
en+fzi2kKyddWoxYiJzxp2oafWc+cvmmKXAQ+9r3M3oNPsMLXX0DqefCt1Iz2EPenpHPutRWegGD
man2Yi/pKmi65smeaW+NIRwtfU7nz6+uqx+3Cj7pPB+YDVHIjgdc7PDZ6YFa5FMDvqsWVJMaCyUB
IU9+rxM3lh3nlfvmozDu+9HLCO+q5+Y5AVwlww99c/+8UfT3pNqRFtg+eXRPvyhLnaYTVRNgtpE5
a/p/Y/vMWi3o3cai9+CT28wZzI7N+GEOnvu7zw1UjHjK/aYBkOD9N0LONrtbn2wxl7ERhdJLPbso
w+9j8l+XKwkfto3sseCvboLzmr641VSL+aNbAQ9Y9Fow8EMcSCclVLNG1MHP0VufU/WmZiZErRdA
N4QYb7jqCXq1gReKJmnfPE9lSGMRL//InOtoa/Rl2Up9DogQslu868pdiqV8Bk8+Ba0ne9k1wFmn
yHY7k+0MmvQQCi+EmmOTs/o34C23H6L6+bYUvAR2hYAl3yrunQAfBZRMmmroDKpGbpaI/VnYadfF
LnvN8B3gZ+CTcQfU/36TfcKD89VEmCnlWiBaSsByYLYhCaj7rV2vE2bWBG/Nk+tAbDbKpXPMjU2P
7BUXcpIA8k7+SWp//XTSueDr6+CmQxV6AZfYMvDdFAh+x3MfDFzgWijqk6DrVB9lfD0oTUB/ot28
bjzP9CZHvkKDITLUw7OjJ928b2OvDfDwFX/XSfAHJx45stFnDOud5jxQvguK5GZuW30CfIvp8R6g
CQqt+8xdnC/M1fl6NDJj6c5bk6iq49cWKwETS+POAtLDGOY+CJCk153K2DgunNoWGRpJhp5cTHa7
GyUZvvgO9uKXqhVbGFSXx0aLe3ciKkFymR0jm9ceYNcHhL5XOfopyMlo5485aAEztnhygYoZPxKs
gRQROa19XBdscnqGZ/r5bYE+sHpDD8M9ctVacOVjMmjDXUNbea4wNSNoRO6k34e8Vt4b458Qs9Rz
7oAfW2UV8cadAN9MvNYARU0KWHpHs9LZOSuUk8pL+hqFPF1xVcJIXFf38Jb7z6s03HJtrDc6xDe6
WiWdqlDPwce621nZJebEe17CDFtz9JY0JMCVlxEcVQJHNmQnD/JmQf68D9S1A0dUCMkZ9ohNaniY
GQ0oiN45XuqvJrWyIVEHcpI+oryXZPd7ITCkinWMVT3GCEikByRH87fW31KASv6Dn16+vCOoYbwp
q9Nedu43V7W0pUyAuIiTXJmcDhIJyOwgN4GbXtUkTQx34Wgi5BnJtnsAi85BkMqrZV7nAs4xrgd1
p7IQti8J2HpGYm+lrziEJHv6tuclTwX7DKprNxHaDYIHxbHV0huiZLUrmkz9TstXGquL3Wau/pAb
VuHHktgnsnbr2OtBNWWfjE13IMweOREizmaZp1+Bs8bTfQWnX644r/+w5N5u/nCeGBbDcgU9m1r0
brRo3Ku9nNdkylOIJDPnsE9MZnfse74mRhUhhh0nEI4v37c7ffsD+rX+5YzQepHX9rNbQN+vtx4C
cPQo/aSKOxfOrc0PmpfLphaxyVnwBmau/l/bYrm2obTfaHJw/IX8xm6FoomYtH5Fj7nrV6n/02Jg
oauMkTeDNVJdkTraTEAPiWkm4zSiBVrIPfpGJY6zM0bxphh8+/3atKiMPf6SOZuUEX+XSsAO/h4z
UyM7bZRmVPBbzfyt2rM1MZzIpSukNYiVZb9miqqYOaEQ+8mNmjVPCKu+VrtQjsseuGKCV+x9PSRu
oE1+qRhOzr/0ck+6IKsXVftLtBT+KJh3y1Lmh4NdhCoIghLZXlea31FjfrtOBZ6YgdaBSnUsf+hs
N7SvKZz+276daj96u6t7TcMDwE4RMEO3VroVsp3oCutUagHSiVPFlUj+c03Op49zDsMgc7fupDrm
JWa1kEEUxnErAMJEl/YdS089KvPyFRFtWj8QvMD97OmA616pnMUejDd/pRGm9Y1CpbsXUhRQyem8
9VS4lGjbeGsqSLsd1RyNbxyVn1EibTud0IoAbudJthbczmB1m6MqpYJkmZZndeZPti8YbZ4ltJA2
edYSOzMHDnlaSALPLQ0sauVVYZB2TKxDHhL+qBRry+BmZ03PuTigweOsg7SGYUYXl6Xwkg6+2Cu5
eb1Ju94Id/IEzJ05K0kZySll4gP4blg/zvB/YCb6Af7TdIc4BLR6zXkBiLCYqV7UuWxMKTVkZ2O6
VnMfVi1dn9QzQxqfMmgQdhUpNlZEYxsDgQDX79eAhSvGVgLUFcxhH5HRZpQkr1IaZl9eqlkmqMas
y+05XRWGVCrzhAw0NUpblwWW/Rkb8HQDY57/+VS+OPud1k4zswoY/tnl9PJTZSY6llrWDarVwnvt
pZstVAmYTAgncC61OffLxIBG6sGLgzkCCKWoddTRwO/Wx2QtOzCr4sA5Mvk5+liMsy0OuCr9Mfr3
ZDRWFZRpKT3Jof+sNMZquS4VyDVLb2zaRlyrZGbD1h9OWldfkTI5+npdu1bGe2ygQ/UCsvaNM4S5
K8NrrLaoNwQi7k5b+CQtSQgRx65wJdK1v45hwciPZTLFkn5ymyNdk0aCtUWPJimD/4suAHOc8Vlm
piw2BjiJFB5sRUJz4BbZ+X26GT4XltV0bhRKnaT3vUdorTXSTVZDIwzB2BwQHvmgtACeP5B+blG7
/2Pw2i6XbwCDY8QofbcPGc8mk7ne7TiCwbdV/j6Vcbb93wUzVBsquIBQ4uylzih2w79Yg8bxiwT7
0+glfWA87bgA2zU0pVc1iVBAYiB5rueSbTMlgF6dXa6V53hcLBFMjnWR+xm+S39IifZVpXkfSbjI
Q5qq3pRz1TeQ2Ms+PmuS10vmv2xa6Cp5UVi5a/jfocjIogRgiBxUqSWK8lvvXalOUnNmZx32zvtQ
YFw6OWVePBYjk4VLhvdFQ0L/Zz8oVBzTU2ebCTM1nskMUfqZgmudLb57PawulWK4P/DBH9rRizW0
hAQZXGHVcb4fJK5K3i6vWga15NnhdZ13ae+b2NzxOTRrLWGrn2dO3ifYZGG0SO8EedgefxbPB1wY
YU1cZNWdTqpoTuOg78nLpIKtXsFhixDELTPsLNPGuwoL+Iv7g+63Sl5MgL4tA4SMHasHMPinIR2V
CRFFqhXKhu+oZLUqq3oosw+tbsD8ZukYFlD/saTTo5FSNXZbd2VGNAdLMKNjVs2N7Et5WSXNdr54
CPrtS7oUc0Eoy532YIzc7T6ElqTxv1nCUk5kPII3bpNGG4/aQc7oKwE++az5b6JTAzwqqg2EANxl
SYaf2iccw277/zKN+zp5zfutzlEiB2KvnSDGN2zE+d7zuj4j72zuiIxyWe+ozn47zQVAQxDLUx47
WZ3EAvckFT4/L+c898ToGNvtnk/jk5y/Qh7dYbjJKNlfA1LYoaP0yKGi5yCLHMn/ISST6OnxVVdT
R4b0qwIwQNs/KgjB3T0EPOt8Z2r2NQsj/hNbTJaLiu0gosyC+wfFmrD2PtzcoSp9jjcI6iO5vGgP
OYCNunSQT28QQzRJ2rjtg1AhZO8HnpjpJNOUFwnv1JzCuYxGoIgHfC+/oL0Jpqmg9C76nLjLm97d
+wKvWQoy3IlJkqJenXL3f4Cc2+lXZ0F1/s3AvGPkPRpom5lxKQinO8VZnwWOOOUhMJNequ5HNEOr
XrHyFdf1+1Crexr2fvURLWab9FgqgvFzGoK/j4HscOZXzKLO7wlCbCsEkry/3Fq6cpaqmwYGKFYT
Z2gIYGMRuU4x8iMoqMhUfYxDA0eCI0XbeX9TyBbLcgSM34sPRJiN5eT+WqzMNFZ+Ppiym1Wo2fU2
bL3oV7I6mAuPbmJ7g4f4VaIF3kWrQ0XWXEUrcfvXmavR+VMDtmmdLJKmsZQzSUlSSYuCi+yqiUlJ
oPvMtFpHdhMKnuZbxHAoPKHOa8O+RkMNsYb7Jd6F1RGcPAderDEgBkFIjOBsiSs+0GdMH8AnPK6+
e/ogpYlABreHJnSO46ozezNGc1bx+XX/tW3k0q32JVUz4i7TfbJsMWhgwGTxWyLowNzAfFuPIf1u
ptwKBOTevND2lVcC4XlH0E12edzeFFofPKRrT/zLf9XKAqK3EvAEtff1nMGzeScj5wdbc6nxl5a0
yMyXzUZMSmY9Tbe/RgiSzDDJrf+haE7tF9hGso+I8OdH1cI07UOcSA+942G+q0m4c/L84KrEuPnP
HMVRBeIVyej84BxVWb021VnlTDjmvG6Lfeqhw9mjz29EhYZ1L2dYydoZZvgPZsLHDn3YAmVFYOOJ
EmLtadxiVU5Wkr/xJeOl2xjlZHqmvBH65djGIb0o9enkXWsmfQvQOfVtgCU2iiVwvFvbKvphZpjG
dq/TUxij6IpUE5/wrOmVf2MIJ32vmfFpRnuypDzp1N8O8TcIvRwz4pfIbawO30M8Q/p9dCCQ8wUn
Kwllejk+sWzTvYqW/UkAFlx5fC0ACCds7WwVHkyI8XUZpBcQWgnlHKQB+YGDb56o/zJ4Z3lz2sj7
WHc9VmqAjm3nWlVAUUlE4+/Vqrk1MChtlYrkRdUZH38PhdTG6N5ZgBhnsG3oLxQ+V2bFD4BNDAZX
x5ut+6MHrmqEZYSEvMSqVwVBA8RaxbaHQJQ+pZ7anGxqaO5H4wUtnPYFEaNAObVZCEKUtzSXlQwb
dnXkWvGdioMHBuuTunZBRjNWddOvXinlMnd/fB4R1hR2eJIhTD/TV/4u3KE19AEUkL2kki1EVnxe
Sgejl9UcivLitM5OHpbMdoNs3GfO68GoP76yQa+ljfnqYRfkxkroFGDONxrYNFl3Xvxpn+Xq9N87
H7Tdeue0WXMxnGANK4YBui10PoS+c4+nH7D6a1QpKOnVkO+doLEBFC8zp3LIrdN3XQvpQIc5fegC
y2VQslLYb0df6BtRMXf5kCc5u2ySsqMVVSHfiUZufg0/w0lEna8UGIuESOe5kLVK/tHA5bEumvE2
Lk+c9vM+JYpIYkOm9R0O4M6Wj3WXbK/PNdG8tsr2UFFLrdq1f7qOygn3f9DH3IejHWkyNZISLgbt
MLJsX77M17qG0OnFTxm6oU7dJ5eemkNlxfMNzw9VA4zRY2iLeuLXRIMRKn0iP++p6ZGxd/+b49Y5
I7fJUOA507g9ZH4xJtT8re5369xixjTuBkHwzVNaRsdhmCMWXfAeSmepELtf5u3NY2LY5KzSnS9i
i3yz2j36xQIS0qWv2q3SV8aRPcrQpPiiZS4tgKJb/n5yVksLpnoJfeIMP2+G/hEAhXb/MgOtozJQ
QaC3JhI36fH4KINSOdSv9rNaXB8QZFaLrz2jf+FjFiMsM/bYm9+V/4nyVKKxlZba/tpLG8Qw4C1/
0Z0N0zXJ89HulvgCCUxb938xR9NVDcjyw4cOJHV3+bdW/WGXxqjghp0vj+sPQ5YsCJQFn4RZixGp
1wAyXCwydtWQkgZ+MqbPYszKiKZ3/Mxi0IEMTerYhyfOriTCDBxeDaVjPUXsHy0nenDdhoNzhPor
UEDEXgpjbFuSJmCGuzah+9RzYdXQKV7GQroBoQzdBQHnG5xUfr/c/k38LLgH389mXQ6102qQ4Tn2
ginMWlCClymE+f4sR+1y+mHlAfMOWgCTJPlkHCxBvO1MZpG13/ZCDgOWENatIqqLwyP3jYicmK+j
EaEQBcgaX+c/Z+4NudgPuV5zBrqhix3LaAh7pXeUcanrrIFap48/d6wxDjqIstkJiVTANDniPU/V
NFtgfurtdK8ZcKMy0Wcy2fV+08Z9BajdH8/hLk1CIWG90BST9oV2AvKBckd5vCyKcQUeL5MfrYhH
mnMriwsz1XW3ryugm8vj8snWGNkNKxzJyBUXWOeLq/KX+CnemI6A9GaomatAAJQIoLPSY7gOlgvw
ZssFvCAdaeXtuvzmoeBbqSGJzMXDLsmJzkJGYFQeBi/OU83izFfzSyvbVlci9ewe5hP/P5IWdUwr
Y5skTgQMPjO1l/OrOLC3WouV+spVGe1RT+XE7lXBebtwxv34JUVBug7KIesDk7uTFaEPMh0p8apX
WLI3wIFxkHWFEd5YgPRy49TX/jrIyvxZNetDSbXGZK14PudMWMoZ8sdrrcuT4ZKO3Pmxi0bC8V5R
ZZIeUqkcXAJgN9j09CFWC4rf73OEXFiIXo6wwkSGvl50g79ZVd5kEDcno3i7DCGgLwajGs29bCxC
g6V4TGgc4GgiUdY06K09vJ5eK/ElzM4s8GaMFGqqGtaZaHnUK6vLO9Knnvfy3K5WaQ3Mj4JUAaws
qq8WKL9es3BWaOg8YTPSfIZ/LtGT694pZ7GuUyBfxH79ohn/qAp8VZ1cwnUHCLez9GpnDKLwLhj8
8vdUasM+G02IJlXNVoxGJOef9Zb73MUosACsUyezbxNDIdQFqbMaLWSUO6SxpFtx6MvwCNsXZL4U
alr8D7/CcsCbqcD241SUrJv/Wqp7fx9wgAXTSmV+i1NNlb7S39YwYnLytItLjnL1QLcf/XA4n6Sf
AlNiuRKlDr5R8N6nfAf6TqbXZyY1Q1WJE6u2sXKS7JNgqGQiFyWhbHaozD6QfJ3QBhzgyfe1TgjL
d4NOIKJMaO0c+b0aaMWUYPYHWHDWPtQpxNuM5nr3wEy17ozmdhRzKqyx8k08OoLklMoXKED0TnyN
GHJPmQ/poAMvoOviK2o2qBOnxZr/OLdZS2sRDElqwOebBtRKSUZR8ztQWRaGVNscuSn2Zdh8po9K
th4IPMy8zqfvZIUDo3SAcLgPQvfAAyhMY24EjG2M7WSyosOVdlAu6dEK3BJAfFSMXAXwOkIUWN5o
V/0NrXBZlo51tNIH/zveriGIns6OKokLjuDXnKJ7OscYwMTh/NtEoT9WFsfq/9R1UC5FDB6PNKBO
6nAkPhWW84JqCOzqjl83EGNGjZw4m2x2LYWl9cZ+ahm3WPU5YHm7il0plDMEMdQTR4Gr3DyDJgQD
84606xT447GX6M298sbciwJGCUKGktKlSAvODc7Q6hruRYK/xaNa1xIi7xSGYgDCnk9Am3BQZspm
1DUI10DE/7mNK54MaEAM/2G0ANSSpvuzVTRFCL0OzmrWj20SBXwyFMn5D6iqscHfxM2yxDA4lsL4
HwCfkhoyK75vagpzZqB+iGa/zVB+Gl2MdETdfS6rI1rh8BL7/7EzpoTvRGZ2Vyv0b5jLHXA16fil
7SXX8QrBjSvIpOcepPmO2azU3gWQbTkkHNDaYJ9uYzGwG6Frwjo5GkoNNIZHhnsQXVDGk4u2I1yr
yY7mNLe6yEL9+P0+umUsKKPemKr/hET8P1YapbfVbvNUbmLiqnkiQkJySZ3da/roFEJ71gEahMCB
wOTSLkoG3o1XMyg5YnBpD2r9VYwVTT2QtgNBusvK+Qn3yZ+dx8jQ+w1NbUm1U1tD/AKWCkchLS+e
PZcnxlLrfO90m+rpmS15f8uwzuPtFbr1SL5ksHo06nsIsry7VSGBbktuon5IVDiFfNFxR+AQYrbX
GWvtZScbCtiEFuAwPl7GGudoj3wuaG3CHAWsHr3xsDXHh0lT+hIOwhEv+7YRRK1TnxnkUFTOUZJ0
iTjiOZedYvapNo3YSVEVfoemzHHCtW5nq8jOmlfhGnnE9g2YI8KXA8lfBOBEfVFVew/rPQ7ovLeE
jIzAa9Obn0AmqrM9d66ilJ8K9MS8BT5R/WJZB0+AxCdisiOFkoKbmIwfVVZISuXnr4YJzaYsRNKg
4f3rh1I7bQtp4Dx7v0zMqeYfzxYi7UtmD4A5yHzP2lWQpEM0+j8o+JLKqSwJfsJUJVk3AFgoFfVW
CO4sMJdDE2nksvHiE/ra5rFDIQ3gjvi1vsFKBz24i6lRKV8DU93AkxspLWmWAuTcEBpyqkVy+wsI
kRcKoxjbmqd/XmqDseWUV9VNUQSzvaeb/9nt1cc8KiRMkNQ+WROSF1AjkKSsDgKsG255Yx3EpO8Z
TfmZjeXRDOM4s9rGJ6Z6xb3L13RaVJjxaNEmrag7QqoyWg77U/vw3fG+Mh5i3DGLM1B6RijRsPhV
NNbEgdG632e8m/hRWvECkj9Xi9LXMto4i+Gn0TRYbmAJMyE1w6HHzlRLO7Wiayt41vcN+RiQdtm3
xVAL5PikEZO/+/CayMDa+tzxbSt4S1mjsRDqDyXrISpBh/lO4x/X97ec/Oir3iWYcp1BEyQLKIg4
X9FPPqsnK1fByqcabwUdY/g5ODsYTA5QsgFj4iaMtO12K5lu+VxQzMiDNadwuwLGWt8ocA0Y9BR9
XY2xEJ4ZbXe8y7DEG27EzOgCUt3i5zWcaoaw9VQNhBAiIdlhKKUnVbpR3lq6nAbXoUQzBn32x4Tp
5A10LAmy6yMT87ScSZrZua1UMu/+MMvpijp61VMvzt+3aF/mdASvYGPcjHoYG+G+Iqgej1BHETfs
+Ci6VxOBIwUOGNLYf+0wkVnnz3jtdE4KLPuSEl2/GndSKes7OnpK2MImzVoNvn7W0etBN6DifUMM
BHIlTASMWMpOd3o83Kt6nZ0aEG8S6oFFvixHHHFqXzl3MBufRAkTfgtPccONcx0rvGp2ntI4nMyy
TCy/j/8L4bGlpQ2TsTuQm6qTIct5YJa87LXGKkdZxwmGfTEh6x9ArU2BjRNxakXiawr/lzpOdlII
8+XqQBwWuL1trICMOVGsi12Ewv7bJGtVFclA+kLjKzadqvWwq3/cXU0cXCvvsIjOwp6u4gIlw9Mu
gaHm5MPhK5GQSuqV8JR31lUin2S1oQpVhQ0aHib6hu9SqSdBzNOS1/vi329CWyoU0n3FODYaC3kq
nAJK0GHzD/Ap1+KvYmUa7UgXtmqVr95l24ctNeTdg9ZYl01J811/dUuEPgnRo96gROOCUJXhhwck
R5HlNhPBuG4ebnNhC9+zeuTa3cql9IE+DnUvlD9rZGUEIuu29f/kT88wyadrpxyf1U5P80NCF5vN
cKBVoknRimDFDCm/iEqwpyhgy6rRSHRbhNrBf2iqpovTfVBBOSmjLF3LRASWMgeQiRGSitOhR0y2
Dvt+wkLmDxxNYPNOZen5oQSmwAU8Y7n0X+Stk0//qeGDAGGXwUq4gNga4NuQAbMa9vxuIh/d3TnX
PLwap5v+CA5GZ3CH2lPXmQSRo5cw8MHVHlJvSHwBVApLsgCMX+gCU80ZdMZoosfDkw4KgKgFy50e
GwV+agi3zoHwbsY++WY2j4rYlHaAMSt6NExunzKgxp8+Xz06GJPwJbmW7k3Prha2QEnO1KKCEeC4
mJMymTq5HDiVjjDuP2j4bM8s/4qeaLqKBItFlfnE8/RyxFRGDy/d/5ebmtMJg9jcu09USivIfTuf
nIpNSLQVr0z9pEjn4ra4/x798DEWA76XnIyVa8tt5a+f0hKQjkKtYcAobL9pHiO4sfs9b5/N9zjR
35EhWuvQjV4Bqpmxb5fWO/Hi8equbS5EEH0L75BP7z6bzrWcnZztA3zBRMhFwi5JGsJv3ykQnBWo
ZUQQMMUZxzq15GeSs8rduZirZ8JOxPv9dbxSbMMmWgMKDlJXooIlmPfOp3SJMpl6XurnWvNzsSjU
y1HdUWyKV7h63PNjw1ewmsG8Y7v6VPEOxc7dSe5LUkTOivgZ1rNMV8BW46jblwH1WtMQrgoMiLO9
5BmpFFHnNU6TIF35olQL6VRtF/OCTZDC6M3A34ud8z3ESSpzQKsojX9s4kUNaKGZI3Nu5eTlT9E3
9c7CWNiFX1+wgS3PU2YTdn8jx1Hhnj6BZGn7iKNggXf4wEDLx7M2PpRZx6yqiphqGj0OZMXLV7t3
MW1R9s/ViiwgyxLR/S7sA363LEQYhCmacyfpM4MqC9vSRr4qd9R3HII+4aIywbLSyb8Z0Zc4LEWt
0EPCc0T9bBiYRvlWfNJH4A5PU/UvUEK5YLQzjCgWdlGTs2PTbJ1JWSI8uExqyUmCrlrmsE62i15O
PPW9+BheHuv/i+D/C4Rubkoy3ulfC9TuzzulKwrXUuY26Hvu/ldQ34a4zPwNSXG+BCGILhlTKunc
+VV9jaMosRcjQxgojeQMoJkTd+N6X0Br6MzofMOs+e4KjLcBB/Ht6nLCL9SLe+9wktDxD0SvGxbV
wVDCzmXBZjMpIw9R3ufbC8VfVlV3szJMzzY9+il4YNdI54Q99mlDw0ER/0Gn1AgEFj9YKt78kJs/
atdlQutu9Tv+mA7tlZqroEQ6E/weDZVRg0Vjy9xx8V8rgXRq7Gph1SjL6L3475sGv7rZHEs+XTP1
YzjRDJALgM9zj1bJTa+HxNEF/D2yie3/2T330zCAC9SZB7H/OOo8ZbPeLfgPw/3fWNhCbcGgnKrJ
9epkJwbSCC8l4cAZN0aKzuQoxENeaWFryIjTOaX4b8TdnsRKVvi2y4VBgqb3OBCp7aFCQ8exHSyP
8RJFt/2HdigOeM8tvleSHOyc5aCl2r5MPjCboFJAX+baBPq1VVMnr6h7jsirvqfoWGQkcfrIWW0u
vKaLoJAalLnYkMzm82M/uMbgdH9pJQ1+3TV4t4CN/XibuvDiso+IlcBqKDaMqzjTJFnMT8ZOTfTG
azyhV8BPxsegXLQlE+uL0u+YZhUUM9bNYTDK81xcFUKN8oRyh9SX0Qbsz5z5fT7cNi3xT7KPlc6C
UJeGAmvs52Jh5wOJt/7qSvLqF8130/R1be9ehAXDIn8znHUjIjvHVGRx+HdQ2/Lncf/BniFJ2CON
8qyeVjce1qtvM+cEL4eBYf1fEhoFqTkW1ZhHQEQm/WTshvCiOMFPjorC0SeSv7cvbjdBaWWj0+gJ
VM9JHh34PV0bhSxiWr13ItvoahozV43mg7ptd7uB1Gq1eDQTsPsLQO7p2uLznvQqW+Q1De+S8XVR
gAr5LrVv+nsOiOpES3dsPNfNYjyS5QOWRqQ0LnknEUswxRx/Q7hKUdH7ACYpWqAdYxYzRDiXBVhU
QldlXjkXTKjnSSY1BGdlpbsoReMnObsw6ruUQWcra+jK+vUQpX41VaetfGrq3I2cmxs1ayc+3uI3
iHfTWWmMEenv54hyFxDkj3pk90yFcxxx6jbPy/2/1lCqA+t6aD9WZWgGTY1pUEtq66FR4OIixzXm
rIYGcA6/0FD85tsYW+0Qso0kP8GcfemPRUbXWWfddWjhPFE7MdqvsbW+gEt7MRT+C4qD1o+KXyos
P0lNJdrCzU/NIo7VTqNNOk68bhzODMCluloqLOdI4Vp/iI7NITJaPy4DX4Csv90Wq5xf1z1wq2mo
coYMyw1OSJouTXZ6dOT21CbXqYM2kbL9vN8wWm6ys05/zrqq/vDDZbSQiIHAu/uovBG/29/L0XLu
gDgBYGto4UPmViI+bAhex77t72fo4UETGJxbI55OSXZRYtUq+JaRu3SCUOepLCsSf3voN96Qe4yF
j9GTUiB74zx4GH1LwRAwNYj8vDG1tECtDfqUuqPllEx7bKDq7T6OAzmQpghRrLvdUjfD6Mznezl4
XkYLNuq922VBCBGZRdxnW2bqxsNdjEaVtMZ/4hPQmzEkxgapTYMSYYLyzWOqHWUhKckWrJeCYFFa
IE59cgxRRoZmw0qAfKndGpH9k9uJ20WHmIRa4jUCzwPs9x8h0D+lBRx2PUic2vPPVEqRDMSux9Br
9+ERkpnHHRdjqlXzkv6YwwodZxmu5zp2Rm9padzY+ymdovcc3fi3eu2WjL3tGue4ZJHUbrs/5PKS
c+R9sfEONzYt5dz4rhXwaPZVZafVYO5vCmvjDyRewGvOb+QmVaaPyUPk8fBhsOFSyEwUP4DZh54G
vkoIJWXk3zQZslzv+shEAdzWJlF1ExY+ZrUeqJIJhS7S/ClntEDlx9wBG7tpMVXReUfIT/vPdtgV
ao/4tp4LstoHJM6mId5OA6oLVT8lcKppSPGCrKxf0ttHooKPgdQ5fjqwInWy2AN3r2zaMiCSQ7DO
dn+9qEyv38IFYenXJdmIvD4W53ZB/AB+1Fqx5jjPn6cfZ/D5YkfBTzpko5y9sC8c7B+6ecwF6e21
hBarey8SkqWMdCYEv2hrHcJnhIkWddDHQCaw0Wi5scpq7UDu4xkzO5GXbTwX+pQbbJQzn2dP8Rb5
hVYRUo5lg+VMzgAXfR8RBL6bqa7jzHDP96FGDftLNmaLeq2KERjRs/vfT/3uTXNYT+gdfvV+j5Vv
U4hkuzh39EyXK2mw3d3mIBulKgMnEWUQof5raooVIT7P35XcG3C/R713cjBT3H5VQnRZu4NEBOoc
+DruAMXY1MZdTqOAXRcxCI3iIMnbrRE1myzu95FYO/u+1edsblHAS+2MnqK4il7fC1DGLmoyZM25
s0JoTv9QKmvaw2uhYZ/GUS+QOqbKR7SPnxmuMqLeF4KjSBXKISQh2nwEdHZszshocIvRtnNMDzl+
tiAAeFWbPxp9qI7Fw7uWUmIXhEl3D1xRKq6/8BP9Uaghr5r1qEiByuIswbxCymnO1mxdu21ERTnL
uhXWHzubn2LdVFm1i/w4SuHOvc8520rKd9Sg27I24DdxTauVbdEn4Ol4kpkXzsBCMMJiCP4760w6
HbpYNx79Jw4pJXOofCKHFb0+yiatZnFrZhvHIHcVhzMnVtNgqqjwKVBnFIzrF3cYynS5Jj3WN7IU
BvclrgoVbo1LfXo6f8i29PQ3t8F0lfB76HJH2Cj6zvxNRwDCoXgKpEyCETQLVthm2rlTgQqkmGTz
S4PHkzn/Vy3LExrt4CPJuhFM9nYoowDhH/Q5XIjBG/7MMHLWIsoQjppc5pzuyZJBAIxUnhH7IQ6x
XMjndzWp1DG9HRvGnONcsJAPSNWUf40gVaTVq1goFRXhnRPvGReFxdmUE7G/2J5hRXBaKup7CeV5
bajcf3qDvuO8XDwytrw76ZfGmobRIC/kGjHe9TbzXtwFwJPbjL//8ya8GLvJ+zpIyds6K17D+mAq
4W2+8PbcSeW2JIad1eEoCD83rESczOZ7l7WG3YW5Jis7L4DJkxiBXhh9CX6gChsFCWLTBHkc5+4i
XOkoT+Db9X/TF9dkBg3WfYal+eejn+CQwOO2FXrTRtFqOz289wdIuPw/DvHdbqPDVJzGs5+ok8jC
6axXQU5KGQoHl0vl0VUrVtNOGGDXg6yjGw/yQVIhDN6rMkPspmta+DZIeljO22T8odZmm005TOFe
5jpXuuiFjSiaTXSrWeEJn8lZigDQmfDhiRm+2cUhQWmPEPezIABqwzc8QkbI50k7yx6U0O30aiPo
xa85sy2+j0QJbQUQXyPYN3HYmH6WUhjka55Z9oOArMfS74BRRyl//SUKY7109+GnwQE0+435ijv0
LcdOsoqrwizU56Ny4pS+Ba08GfCpW2rEIz5wSScVjiYESnqsOhERjT75L8JjUBHAkmnHHbP5tcjY
m7DHQpFQDpkc+Y4SuTVK8et2FRi8AsUFYiPPddpYCXjSpR7JpSVS4Ikc2i2JJNz8Q5XioDoez/1P
v3j73vIM2eA4l59lGZ5ss6TErGQ4TVUOHvo8XhfeYYSp3OkAE+DcGuYFTS9bq4vXghOcId0geOuz
WFKe11sZsmXiR3M9HEhKIh8DJ9Nw4uDv/69nKV2z6kBqxA5y5EeVxq8aw9WB7JUNByA+Po99lyyB
XdeMEuYvq/nbZrDrnPlAQvDnZzPfaEQUt2o+k7WZxPIhZ+Wmg+oHKtlI1gYW5OhGtTwxmKnbDSSm
jwo+SFiZRqwUqK1xt+9rAoOqTQKNUsHaN2/lF6R+DesuT3XAI4D1p1LWDTWdgq/6c5+VkmKmZVHj
U0cBSv2Vwzi83goMa13FkVVxbzt7wkoH3tm+rzlbomDeimmq88Fo6vD2M0cYvtTbm4LLZk9q3SPv
lJm5Jhn0qcgCeShs38fDLp805LJBMsVgWtqN1lvEav3ozaMZEMN4Zk030u2WnplTdEKoZlCoMctS
W0Z5e0TeSXY8VhMYaMCh30yB6diYnrRj5F8vGWF8CabsnpUj/0T6iCbPHLPa+eN3LYd+Tz8gXOCQ
EVxf2a+7M7TK49gUuoj27cAO8fV8uo18wtivK+x6KY8Gec+u5yQDcuFY0sArzVeBlS+uqRMDIh0y
iXmJZeELnmADiRBf/ZzWE4deSXyei6oOXcdkAPdCgHb0p+jq7yNfGqq16REBP5WjOqCnBlzBKXg3
/D+KbJI7MDZeVzG7v4/PTPNDPHkZd5r1/NSj65CORGRGRbFCoPHLVcOULSy/t4iGTloD5NkeaKu3
0TevM7Y45AxtRKsBFNXCgiFlCuAXW+m5gUdXSKfbpr1WCc/I9Drh4kigA6fhJmhBc69ehjhpgQzG
k3oPWW2wLErbKTVlTFY6W17oTdBWvXfBIBYhva91D7k1B/51cXgROnOVMZJNN3SLJnpzzC/ae+/b
2kt9LpbY5rkjNOcc2XOhlmbWNb8N03xBYqp4XrZ5XF3u8I1OwaXqsmGSzFL6G1hoqIzz+Z+iZ3Ja
kj+/9/rzwftuRFDoT/YiMcuYohSsXFpYpjMR6pHifWO7gP9sbpBfGWImzffI+xXt3LXUdqCHnzEG
AXhfg0yQZ34X37m8OJwW0LUk3fXcbrmKGumNt+ExRwhpxKT3a9HCAdWkwGO13OlbdzW8xZ1Kkh/3
KmizdqyHR+xrY0hgMn0GTC1RAzvt3zrW5mFw8oj863IjdBpMOtYE21iwguN94gDZuutztG2jzqpV
UpZ1AsJfsCLm/WW56zt4umOmoddOAM5UQ6qxUMei6+Rt63EQlqu8he4spmWptGLEkDW5WrYnhtve
UTZbpfAbLiDsPEOpgD/Sr63j9Hi8pxIG/8NSJP7Eza0ukMCbzPVsIoU9MRWnQEwv/Tsd6IKOKndL
DYAfRirfI4TPuDHo3YphlpG8Zxgut4i9a5SSWR1n0wemissDmCm+vr38Ly2abSUgv71nhzCY4IVU
Ifb4qzUX4UU1LS1j1NEkj6Uv0nDd46YzJIN94tCrYVWfDl4npLhyNR8fsAsSsbuTS6bZeyfbMjyM
ZOvV1G3nTFrh5mhq8so1nyPNzr0pXeFYMu/iw7Q4/qHIGLfGiPsaoC/se0kPRg+YoLdlHmzWp2P2
0g5TO+oM0iqBUULo1QjhDsS2SXpK1mSRr6FkvV0Iul7CNZtvGuYxK9PFJpmpTy7mwT5Fg6l3oANa
qrHgbF/ii50GLohoq79llCgoU/DYEYQjdjaKaF2NMlko7CMUIoY2596c8qkjlaJGHxRGpyY5tpiD
3lA+q3oXUHQe4J7U7uNk/PusmLUfC3KuyI5Q0PfVr95Or7/zvclmJC1RACm/EEDpPKcz57/IF/jy
op4fAdgLTTmyrzt5nY2kNiIGyZ7D6EB9x+m4Xeb9Yzr9XjvDndPJFBkvMbhZMiu5U8pfBF4vpTNn
mNZWfRQu4ThC2HNalanW6uQq+Ykl4a4RtwQt6hby40MNzNqn3WhJTfRZfD3Rexjv+CBN9w9UMGIY
eJUK/RukkSs7E1j2Nrl53wfCSlF1C4Qn6bu+qfeQLqanSGQixlixzpEPTdK5tveNekRV3yPDdPSl
vkY8boXCLct2Jl7xwSVQgwKJ+z60HK7nwT02FxIJXGW3DL39AgPCEWh5CxOPH+HRhPy6reKUREtk
DrlP9A7S5DLf825k6rY/okg9w35xYCNPhjqV/28npQf6DIT4GVbvT0Txv8DR+/4+jW6Ve8cM0acS
vWZyXmgcJsb4CYUIPGedWaxaieJuw4hBcPJd1FGMeidS+8/JoimAB7ERTwtl4A9AY60r5aSR2Z4G
kGHXEQg1LoX4mA7ZGFcB+R8Gm7cY1u4ZAqoarCN/2ASBgRzS/rpDbVds/HZ1qHWuPM7E/fFB6EID
5ePdvPcnEK19mfB5c5ZvcyC24+JU6x8d9DUYjTZCjGgwwc3FdeLzqKRjL6SqsHsRiyyyQU0h5Tnn
SZpLgez1Mp9gfN/LT+ky64npiKs+ZDQ2JofniGoaAhlw1YAlSIdOGAPufKYog0LNwTUM6M1r9OBn
i0Xq7lhszuNGudKxwF3hHU4wDbgZatqkFlQra/ZId1W0+cN1GKaUM5HUq5UqYBZlF7K8u1THIHto
m4YHmqv8hFHn/mUzAiZIK9+weaagfmW8F+46SdRAH5C1CNX6Ed8ZZbUYAzrl6mNM/Xdhe+EtfgHE
Ng/B0Zc+v4cux7gmvyBFGfofYnM3/7Hq91MYl/fsxyBqRo9bf9jHzkyAFGfLS4B/WbMI4cJmyNT6
rqBZyGuWT5J0LONxMhrddfz9dFzgSQ/0+g8WZcT+bCGi3dhjkS4phw5vXJrHMr28gV5XBAZvsC0H
GujOueSE7auuJHCGFVUIJ5Cv0nOngSU066FfcHOEC0CgF4oKdPHUDwMUQYXI1ctRQyaJr86njo3u
uSmA62XEtxXXl5Ej+2Z59e+Uhr02SPqXsthhP+vMo3FKq6s+80SqX6j3O6+mEDudKK/9XYtt18y1
9TtTVTUrD3MY/xStLMbM+8YO/aOZz3zAuBANW/Xb2Iss6vfoPZHpPVOL17xaVaDelQehtGM7vP+h
yjTplfoDZEkRLR/Ko3/r6PlE8mvekzpCmpcfM7WoKEBQzTOpwk/ONvT1Bc42EwRJvp/2JPzxUT6O
RrSpNYIFbIo4ax/oyurIT6r+ufViUmc8a1/DOoz9WSyh+JqtnBpxIrFbgOQ04LVRl++RNllaBcAs
SnXLT5ulcDEWNutmDTIIIBK2AjXtgIBYWndCdT81PByL/e2CJSHxdHQne3zHqL642lc1zbj1pnp6
nTp1KxUV2cudvCbzji8LuX/X+YEPcDyu83h5g18Fxco8VI7PXFqzweXn8bGV5NB4uPFPMJ2wE+sq
caWFr7/TtqBkRVVKStsItepMNIexGi0UT+ILFGeye38hWELbmbTRzA7oH8dFsTqU+bNj1iMmOsRg
X7vVkv4HXAGfh70oM5RqSkc5hizRvavXpMyaIK6f9gfytsHN06AIdIPNwGAsnm+Y/NC+VD+b91qu
fcjmJkq2VTtIykh4rLAZi52zuHfi5Tz9nht9xK3mC3px4at02y/FiiK35AzOxTZGtE5eTe5oa2WU
sgB8+RbzZUB3MVhsMKiIE3u8gOmbHZZVkqz8NH0TIWTRRNKcUtxLyRS100lhIcuemytslLIIvYHH
XZwsFl9iTKNea8dqV60LduViDV9RtbhITELwC2eq/sv6CLe94n5I+i0IbpLulvych2A3iRaJRWT3
Otf/oEfmOnyOZa+F81WZWsLH00azqdWXo/v52Aafb69dmVViS7NAKUx5LpR/OYZmWDsB7NnsSOyv
sYt2AdW3Y2/tT0IK3FRoJ0+xz854NppTTgNNmkBF2LnN1aRMt+xQKm9iigGE/SAdmxZkbm+slYkH
EuQqJaggWfrrXA+Q5w87Hj4Ps6+V6s3xSwIbh0eL22n2AtKb0zHvIn85JmvQKOgFkKWKBAGGXtOr
IsU7viW85v0itgh1R5zuoL5Qe9vQq3/1qerFhPlnExpKnkPYjMW7q7M4JJnr260e0fikhOxW0Pkm
89eZ/welMXV2XuFxiyWQfFZaEqcHDJfpmiLSGxGI36Rmp/p4SxQ75SN48Vih6czFkSvzm1Hcm5n5
zvIBTaljdVRcsGG3/5hWMkErLvL68SjvcTfxQyor9ptyllJJ7zomNLvSLSWQJ5ZLoC8WJJsFJq8L
Ka7Xwf4LADzBURcb83ohBnnhELLpIBQ3F9iwxLavi6pa7UsFAGjHMFyBabUE1QzPPZ0qFqUv6f8N
g9URoI4mYqs1/GUw46kOPF6puxCGvvxB9nWNujaCdTbQ0PKAP8oEbWm6AwjJgralJW/jvYrwpA8d
c4pIAX1ospPTgAoYVGJ38momS7hHC+KdANsQ+f+J+4vM0khrH8btouhlaPuXHFCCc8dmRdkFCsir
EQ27Tw2pqDeIs8Nu4b8o+ccQ8zxIDDwxaIq4cq+xk1rOPtPr3tVR9OxOpnTUeSuGd9K9lTBlOWch
NdxpDvKLbBMSC2mFkWo9THyc/HIZHEVH2Qi7AnA5P6YcLbo4HIauFraCiShHyYjjEKJ9P2QvH1E4
bvryUrKXsZgXIH4yPMGvkuFYmmnLHj6rrnrZGcyXELOQ3jyOGQbuBs4Fnva4KhBexTV9pYtqKsKW
YSaKhzVpRNYArCYDcQ3LTf7/uOgyZ73sODNbhDXgvMNwGSk/tlmOzGU6A9wRr0dWrq636s1Ba5BY
fOvcL7lqattjfJZApxwTeyWUjjvdzE/bvNfw0n1VgmtVKrphGiH5zY4odoCDKKh8kU8JlqzlWAV4
an36x4cfswew9MMWqZXmGRBT9ab9wCEA9OYLMAeBQnSl4XKAzMIhTm07LTuSu3I0vCOg2vSM3a6j
CNluuV5abDILasR2l59F0/0hxOr22RUI3KxVZ5gj0Uaql65KBQFqpmzBWYgjuLZLciH9CMysAwOS
+hE3vgM4jmcEa0JoerL1brHv6l7oOWPNzom09zDwgB4E79MmHqZ5R6c6J5n3zhx/5ptHyxw0cimi
AsiWlqIm43JtpVPstzIsol2l1K0R1Lg8G2zBjmZYiH+h+pDHO5lOmMzTF9VpWRL9/n8f+x27d9jb
qi8k4siwNuSzrSaanoEaSZoYEsON1e2Pe8V3yihfZJA3KilpE32C9Cz3LtxGX0/wgwFjg+xbI4xy
7o9X+x1FN4lc0bCJzbRt2uS4+s0Dx6kzq2RMSNLgGtu8vrcMFRRtrxlOG1JK4p2ImgWT2SIE578i
eR41vwF5umYWWeZDnWSwKVzvIjjTwBWqO9sxY3HpY7yYBTe4QjfZaGxImvljGU3sErWUWN/cbS1E
I6DkkL6mTgcM40pJGjYEja1KffR49bHj8T4LGgzipVSGQsvgBq3kPPeCJ9Nr7e+exK6GhMzkpJEP
biUji/5jhAWYsKIq6j6yjJMFhNdG3MEXI0CIJxJxY0a1d5HSNArbXm4M8Eoc9JYt18AB9W9NSLvp
PW3XfN7hJiq5P4uEjNwV6mys/7bAF2ACJ+N9aSaRNvnEDHQK9CS4iq0Rr0k4jC94fwy5PRrTUKoY
RlGZtZyNF36tU/UZHEeNxKmoj6PsOA5KBbzR1daLhDbNtyUEWWvAGcSqTOwX8F83yhm6p4ra5M+Y
OHxuk0+yaHIEOERe+YqQwX9NVvdP6GLDQskuaCcBatjYv47lDNp5MyrlHsbd/QLIm3QVTSAQ+Tfs
ShpsO1UJdUfoejQXqL63bv041W6iuyn743XbNTjNR0iCOrAAplkifhkrQ6gYt65biiHPY0zOmWtn
G7XKLwZwWmQz6FPjE9ebRUBWt1bgOLqaoIuz2Cgn4rzUBnX7M9CF9B37jOAof5L/XO9EDwixc4KV
KOX3m1t/5JMuWXZ7WwnVc2feCaqOGNROPz8bQOood5UPrjdXyAxozZCNDJ1cWJyHjVOh1eLp0YdP
GaneJiGCDx8aj9D2ZIzf6AU/TYGAbCk1lg/S3ovYeIgQqsufY7LRTLcAuxArKl2h1UWYBstOCUsm
JDotqik64jiMI5ua957HSBK9DW+NWLJzPsPct+A1Oiun9HoQP5EdzgyydkFpbs9XgrBh1nhw/9gf
D31913ewE+noboZngVjAnT3aKhHtm45QKyxd8bV0/DnRGiGJZa0X2BaizNfy2EDRCdwU8lYjzPa/
L6kmBFtce/KeUqb0CJ3QpypcOm5fQTU/ulKvp2svHVMvLCN+TUS9AvlDL6LBwqOOvJJ1e3fP1n9E
edJMmqK/yCM4DaYKv+oxO1f5blkMe2W0uD5ahhqvis1VMeS+61Rz/nkN23MvU9/PY5IrEWRImUZx
IKDb0hAT/ZE3LzKNKYakb4wuP28m0IfkEpmWTPqgamTWApvM+FlWXR+h+uklyLfOUB2GKDvaG1J7
Fz/KrUwWa/pbhQRE4zKflI2kxeo8QQ/SZXlrTDf79fKUBPR0joCvtrmNhV5jC8Pp7XPjalqanOfW
oXDSrlGz65o1naANzSpIFVONpBbrJupEzmzvmq/a5bCohjFeYHmE8+LZbwjngN+57QzP/cTdEDhx
GzjA6zHXxyE0mypkwh6u3SVNFKrIb/QhVMhGWmAkXI26/4ng/6uo7Q4wbXFh9zfQ71t1Cm2YEpBn
ZSXyMOJrUNbdg0iWbqSNHu9Ne/499Xj3Sk9LCVEWde7bJj+JOPH8zcKmDWo031RFhoxdU+YJa+V4
HE2ZgnCax26BA9BYHdtowlYqRAk2FnGZxcLc7y77jei5HkSnlyvU9fjvAB9l0pdcyHK96m4W6QSA
BVeKoU+Bc74YSB8dUJcJB7jWUPdqTVv5MPDDo1j+wPvOHn4bmIMUYxLC26jpYQUTn9xL4rYoFRHO
aLxDflzgX1vvuhcd89jLxmc7Q4RrXSsKlFu7Ird1QF2iQqzQckKcsbDqfutfRvcwmv4FB2i4joor
/ZDbCDdG1S7DGuLAtzoMQYa6gcfdsII8225B1vznBX9HeIlYREQP/tX4HYTVwqdN3nl1Wbs1+0lj
O+Ii31XZVS4Wyc4FaMySnKff8DeuFkmjCKCtQDQBzQGIPUsgha7XMqvLO9keZvL5UIDUbh89kCL5
O7Ngy2rGGUFDUtVGRG9wcPeIkOB9qod5MHR9VCCvCNf6ihlbKXK+aWOhtY0vw+xg9OXup0V9mXuF
TM0Ce9rSeWxeCJ1S1hRL6uKnjARRGZooo7p+/TC2HeiRzdjVRFKazlmTJGoau3gRMzCcvbebIpRM
FgLHhwBX+2X2KPz5fJOklRmLEan39i9uNwGRG73b4YnAjvSdrBTLq09qrPJQeHwEn1EIhxQdYrEu
9GxGkfGf1dqWuonCEx3s4Oq3y+NwjURFXaIMhReM60OYcB2QOtjyR99IEEH/Zb9oIJuYY+vd2fDJ
HL/38S7moWh7q/zwYmyuiEw92t1CbO0HCdOwEv2OaOo3ytL39zbi5Gxnl746LHSKI1kCsv6fw9I/
pG3u1zNsVUJI4GYfwFpiVNqDLEJrXuzOL7wRTJgdtDwA7Dhb7EekPyotPxhgzPWrqDkhXvv2ZMYO
xCOlIKbdTpWQtDPB7y236WXDo1DlRvylx8y2GdejVHbMQVmYsE79QdbJznUj+TmGfozsgdWYpTZs
K09hj0p5Qf61YSygaMDPfYTs8zUJ3tywa7FdgDfQJ+ZhDTdvaHaBbMI/yhiCbKlVQyvhAttX22ub
DQuC/7v+qkHCjQHx4q+z2fag1o/wHcURdXV0Wnfd/PpZAc3AgiB6p3GUxma/23VUdTqUtbXY4ruf
BABlVqaTh9uxbYNu02WivVV61O/jFE9VZ93B1pYPM12FaIzMp04Hg+nMXCSfQZ5bJAmZMV6OLXdz
8DBZZemM6Anarolyh1N5bECRydqpDaMeCUlQWQe4Y+wNQj7gXesCW7e68xrYkG+/zkuAeoXQz/98
5JBiFrLBb+IcHGWFZfvlyHnvn6C520mzKsyeDNSra4fAaDrPRGPYgzdjJKxhUT5lkGSbCyxP1inH
nzXAvjg+YLBRdyDfCv6w2MtriSnv+VHb6DZHhGwnANIR/TPDS60rIoEWU0v275EYT6VpyT9rXwQK
ddE1UZgZSmPniV7Swd8T2Qbh41eVLMYkzJO4wzFV4bxFfs/MwaJUOxmfDOqhSJgSF/T36PGxZQdW
fT66IQf5B1BAzr0vjzlFoSa/7xjSiSQ3q/ZKjLEnAl/7OmqnKpxNpCKNdFZF0zq4p/55aAuhuhHC
z8e294KCsuQQDuAxRcLezQZPBa7ig4A7Wvg51PYDmhBu+r9bFFjR9EKz+u2mhJVD2y2OdDcm6AJO
d22OQJASlUxm9ee1+qH+bt0YGLtwUyS4//Dp2n8ESrAOuwRpQ/WK4mYFYzLI7r2lJarn4CHuw1CX
cDjohc1drXqv8QOpq2ANkUjdNoH/0YJnoCUkEDkJ6JHvjmnXeVRZWB6vTKXEpuEXLmur3IOW3xdy
Pmiov0yS11zBKMsNS2g4iwgcw8TcFG+b4S2/XrV7odcz0oRBzKIqhrepbx2H/E1TWZ7YO1YB5NqW
rPL9GmsKUxQFOiMrWKa4mZG9+/IYTW/jwyA9W4On+ufJbyKVyg66x2ms1USK0m1SYsmRwv+4dL82
mJ0VKKlMX/NEW7UMXFvOXztpjOk+t2dg5l4fVBJN7v/cRnonRqBbvXucZMP0aMxOOkItXkFPSdQl
HTJ+r+65rfbNN4wJ+Rq0VheiM8a9y35H1ixTUWnbpZTigTU0yIei3T9xGr0urflp49XVv1Qgwwug
qa5HJBCWeBV2glLIeUl8Wy8WBwO4ry3Z7EBu9kxQA8RJtJMmSniQErHUj0qyIZBKjnmiOtD5Iv5D
eGugHKuIh+RJf1SLyaKVtiM5pZlka/WLzwIzznTo6K7P0Mdsam+z8vrWhZbE6i3qSRPYpFSjFUbS
nugV5m4yg1692dm1rtNRcz283lGVkqHLdVqr/2+1W77ULgkS6EwNOpYRl+xUtBPVDg/PgANFlke7
NY6ZYrpe0myzLxR5638Pp6V0RGeOwxJbQMi5LaOOp6mlByI5MHxt/acFpsre3l+q7TI5HGDPymeQ
mJgubvl14pWoyI0gkKFI0kA+QZ4qGUEoSXbosArSjVF63pTklO5PL66S6vVNqizbNcazTBc3C4ra
VgnqUtCdxsp7oTHwewL8yfaoZgSRGodBnr54uk9pl0XW+l6FhP8QVEnYZ+oWjuTMlC/YtsH1eyyF
CuTJtv7Hf0wvFMHLgGsDpkil6oLLSWBsvoDEMGBSyrLMu6aM8vv2SXi1FgKJCBIJPjMTevE7HW5X
d0sgbk7qSWnyVSznht8lPboz5EfZKd3eb2YqUCPfBb3SzWqvWfSXKLx/FO/OXdVbZv4kyeK3N3jR
OA5SU6YgWIPqPRvFnTELoG92prkyDIojrisDwfHdVuly9ydG95BiNXKWjkhkOWhq3rqewH/PD6PO
oVhrOXXbmNYLyAbkgPTnLf1lglY10TNFq0qyNJ7lo4aWuP3C0NgEdxJkubBlvWuzlJz3u3nIeXlv
ufHBQe8u3ZC3GgQhZ3TwVzevFOOs9nk6COjG5gU0vYLEioc81msTXy5WajX88eUNdgtTBS6aY5p6
XdWMbvteT7vVhtPbb7FTWCSyfSUhCZKf9ZdXCamNuRvhF7XBrFen6nEo2sf8iXisRNXqBGuJcbNa
lSbAAy4ctXQPsYRqgc/gI9K2Tkm3MEjgWNUT/YpU83of80tMIlJ/EgCGdV23SdMb6k+QI6/KS0IV
JW3JJwpnmMjqFDnovfyMmV+XcTdWRI7BC24FnbzLKbtU1ECPnXHM+hvnLst9ZJdtCHmwvsnSNSUB
KP9aiTzWxtplozk58Mfa2nblIGfz4oOPPZ7W74/Nohe9/dtKABXzN06e8dsWsd1nGEUuJhLS6MdC
ns0rOn5MooUATF8aJ8dkFOCoNl7zfupiS3mIyPZq8nvVyYL7xdeqLCWbHLkfuT5+rYkINW4MAGMH
Hvm0vrjxUFItR8wyL2AX4sz4q9FPBI7c6Mf8fx4esMUEdb6qPpPnOxF/4Y56bfnbYji8casFGSm+
MoFn211rGpS8rLcv+9UHs2EIZDW29GJonUdV3DMTE8zj6i+d9BLmEKAHXGmXRekrm2Eri4lq/IHh
lE8q78HpErlu75PsgjnmHNWWPOVLqP7V9NY0gcPVqgyEFSB8QNUfbBSIA0kJGLWm534qr5mE9b4l
xdeHT1lyO07/3lyzy/a1TQpdRIB3vNaectyScpaRyjD5Jb195QSI7s+WVl2JnQuUKzUM1uMCbdGp
Z/OxHPeDThYfKKOLwB5f0aC65MFFfTg3I1Be8YxKEXxQ9ikp7m64gTUY2HIy6j5IxOtqUNrg43ad
mVakqQe/sqzvluy1sFUwk3J4RyG3Dur7nVt8QYAi3862vG2KJI+ZUOAikB4HTPUPt8hbr06xH5ke
F5JOJqz+JUYQEmXR+6P4YNUTxs7AiBIViMENqx7M+8qjdmOaiAhv8VMOfo+ejW6LQ63O8a6xcFnz
mzdWxbssGW2hrSKd6B0afK2iCsdWvV5PQ1+W7f0CNFix9j1Dcz+IJq6tFjVfBtDwdW5R1YZlf8qh
XMLxZXnyPE4d0ohvqo1SFUWhTC4bOG9c6xsXWxZCCd0RT9/p4se31F5Vq5lq/o+IKeZJ6FXmiRze
WfziPEpuFWVwcK4nb/jTfAuftdSnS5GAIC7ogpfhL+R8gawAc32925EXpxRqHO2LvF/8FD6GBySt
8uUyWmDoW+j8XPCMmizr0qQ89yTi5o0w6Nbpua2V6OdGTCpww0WLZhXsI3drzrDLa52jfyozD0SD
6UWoVMaMISWZVy8nM76uxiQHVGlAp44/YEGvJ9RvomMbGrDaDvfWtU3ckJvMbdjnud93xuTcjaHr
LQqMIbT6+1+h1VathYmGQqskpfm1BQWL7vgJEJf2PUPvzmk26mXOMKn9Vb2eQWbbwZhgQkVVj19w
P94dF17Txj3B7mBUYndY7ia2HzB6JDNSPtpwidUGPdbFnSxQIXrKvv8oOM87dZjCvXCnxrvwAaoF
e2tGCINP8kp9eGnZrORM6Izl6eCuwqtV/DdvtNF8d+oDnDyreE4aii/EAXbdRmLFEFUO8y4ArjrN
RMMZfrk8g6aAUYIKH5XOEkcwcZOIBN1dvnQIxrDMFUDtBqc3njrzAexf6Vt76vuSaR5CuR3AmtTr
+toB2bRyDZtB9eeVp+bPlCWDwpKlrfX5myHGyZ516JUXXZEDO4ZxN7CrVUMxqymnjqi2LV/n+7G3
AjUij93i+CZ5KZa4DYlzE+fc2R7bQIi1pP688ow7LWBW3EcMuLOhrEJPIn5C7d5xVvoM/YFW3FWu
LlXzlNb92chwK+ondPsn7mpmdo8e2ILVpdd0dhOHPdVgGo0kyjDdhG50INvG6OuuOsI8dAj61Zn0
D6pyN8ZYiYE1RMwE/09ptP9Q65c8UhsmZK+Gfm+pgjkNpvJ82atOfHetWJoqQouRpvBtpTRw9LII
HIm19HnBKV76GsAQAr+ZtFizqY/xP31AV+JgMPyFirfAsmcfhiZ0i0H3A9mgUIpx4XV3xRfZZK/O
aHtYe2OCCidmzQY6nXznswLK7rMTqEogAhVMrV+cSqrpwBICJmC407lExIg//5fcrStv13ViPqli
t23WXmrfmo/geAKd2lMrL0f+gzosFPl5MwokwkNwN4Er1fMqkTTyTO6g8ZjzR/L176BSf6eMXRp5
ZB2p0g8D5qhZUXWTDB9CJeVcW2aqPgXg6e5t7L/yV5CKhG9mn3f7eW733AReRKdi8rEFxplpxbgf
bm6+8CURRKHLzY0LnDOkrohIR/OOc32mAe5cdV0zLQ8oMyWy6k+gy9bN7QGjNRZXfaajSVMSS8Nm
Vfg0AKTISvcH7aO2fFbuKaOmi461ricTAe23C34VkSTJruenbEEXQR73mzAuQIy9VpsCitbLXMfx
L/RjNu3ZN/9ufBB5gY94+RG1kMnw6YOBxpsv4ROzkhRjx2zq9gtdOD3Hk+tcoOIQp5rmYy0Q1un7
XkhVfzZU7OBaemb5UuRQMZAit/EIUdlBRLKGJ1Px3YqmkXwt5xFVS64YVFN1CSrhdZ8+S50dQhB/
Kte3id8jGEL/y/AEEq9KBrmUncWUCUrUoYv6mXdCRIyPgVTfezHEcqIqxfmBTFa1I7SeN6+wNke0
12BRW2quNDRn4bG3KaZHK2IpfjXcgPrexolw8z1GaGnl2sMcuPRAjEGk2yxw8U5XZJAjc/nuh6OK
5KfPC9BwJlnlcj+Y3t9CWC7uRrmxYRmypH8kmIwnvX09TzjF7F59Fc4VrQF6sbBZJ25XWfnLQygD
yidNobko2fbLzfvS9lF8agKj4ISn3jUTvlj9GI7A7Ot2iK/JzsFbYEI3e9CYN4rNEklgLK/TWT/B
yy7H/b2p9NeBR+aUBOuaKvjl9ciDK07+LNj76AdWghfZyp9d3TijyENjvKUUkadUoIbc7gc4Xu9P
aS6wX9gAX38xq4a6wylDNQCKrnDtd1sOuJl/MUsDMh3BKbGK33G+UCgV4hG6dAQ8Zyg4FqK+Vu5e
i0brDIKXSykinwp4kO1SAX5T9/RuxmGV2NW/aeOE1zuTfsZCn53T5/JnPqgsiB+sslPfePi9BHnO
sn0DZXJ0x9gjx9pHIeYT+5qEq0OC5PodUImc9+ocYRFVpvEHJEXT3IqU5g7EdDUHSHEEKkHcULXE
NL+4XWO2E+SKZwrT7iGBOjU4Z7XuENG8eoYpykXCrT9eM1ygp6/StiirB4cpQ41QuSrSoSd4YEZJ
LEDRlqfsBzYZcvAnam4rlQTW1U3T3Gk+dhYEnEuslHk774CcNN32+7IIV/SG0fWjMfc2G4qA3/VG
q7xOKHSrli3+LrLxDw5pyTDoMMl4+LejQbQONqfoWWOjWFtRzglrImRVkrAFunhimmv8POBtls4x
bXCLzE3/NZhGhlBLnLdYPyaqlCW2jqumfS2nDWkEAam8zX7yziCDieTYWLi/5okyZUOC5C3O4mtj
ESgfh9KY0gZhbU8LjVTqQClejnZ6N2SxxSglChRmTyo9qAc952Kal59l5c2dB81KdQDeDfz92506
RggxDUOGR8usPWLRg4Ij69mD1U5IvWwyiJa5D1uZAI0aVH7Nf9DGlH1lJlcUY4njGB9hFQ/Tjzdm
GkH/C5a3Wt3cjyYxZJuqU/cj3eNkrVrXNhoiYcT62jY8sx1NppK9MFwKnFzJRNjsE4f5SSGjo2rs
DeT8lCt0NR16nMw7zLrJWaXDPoLRycz2PRxtZE/536jIW9gXTQ9s6EEmNhX5E/C8rWWPcvd9qyCG
XAEAlfOY45aQV4C9BVt82yYfmWCI3Opd1aOgExtiO4HzYCVE1AVG3tf9VXhOBboHJzn9K61JyKdM
wEG7SHfWV7L3/tAIbBgPyoXD2lUhm7KUHg9hlNbP57QBZ9SQu9Tmq75HmeOh5tMs12cfMHILhdya
rQkc1PyVbMtYLTWHpstvTWpkQEdRWnGPDxwGdPVzDsbjywUAklJyJpdE17E3CQ5ybA27w8qRltL1
rusNbumdPPukR2Lm3xRjiKZncvKX1sTbF7uXKeXv9jQ8rDm7QAKYrfxwxrz1LHBl4XHVH8K9kdgB
pz8hQtno4aFI2nE+6LzT00p+opUDZ1msSj4tBfGPoWt9uJrN8GP9rJpdGSNk6F+6lmvVsT8Lm2GX
84nayExC4myhUqLSnLu1EZbrfwlliN8h/eHhikRy6YxVEYbv2IGohUBcGnRkHKEU9MaKymaaazt8
SGRWJB43OG+pljwIZaBA9b6cl3/fjVt+ZbFlv0SvfjyYKHp6TcGSgmzA3psmA7nKb/q5Pm3GEG/7
k0zqYRV2l3m3eBolA6ogzv7x6UUeECT0jnjbQHa0sglRz56n3gLdHxcdu4+bAscMAp1RU0JyHNqD
38iNSz0YfeysefDrabmXhT3tmGZAwD4e6tN1MvuUOdqXhdlSMLVyXXulaRxIjaYk3Xfmyr9lPy+v
3FN2R687psHOv50n9m6Gn6e79eYjNOqySBP9gjBOfSPng+Q8k48RXKNrdm1QO8UWtzyzo7q1v+6K
f+j0I02P7yfDyZ/n0/yeFDeGyIQ/HiVq8hn5h+SRYWYLT3dIJxAEArnhaINMSfRLZgGrxHSK07qO
q0KOQccXc8J9RPO8x8HiFiUoMbvQUsNxj2O7UpIINH1CmA8DFNBXCKzMrGpIvsEe29JlJLa7VJLn
CNfhlfEq+5uSYO07bJK39J6hP0ubUibqYT4bKd7Vt8vNPrIXPvO/3zO2/fppFQwjeGoVJ4phhpxz
yaNRwui8k0kBwVxbgj3SgCsfhAHifdrJ458rGWS6HUCct3J4tGYoImeZCS3j6w7Vu9YKeByJPXwM
vM/dEuAuLaYigV/zsGRZbjqiY5zOdLLXtlKaSZctfEJPVbsz4hGXwdWXI6s+3d/QDe8oDQX4W+SY
k5QRyRxdW27fzRzoSry24Jm+lLqAgbs2H5ElitV9uVjO/kE+/KlM29xa4nfvE2tx4zZkCUWQ34bp
Yu4WKCdRyXx1vvSBCEAVGv/GH0plz+P8xpXAlXzL/9ujok9g0fHf23WfBAEcjjjqLmPA1cG1dPG8
FRr2uUW4h4DG5I08jP+nRcp39tb5rfJyfzRQvx96qsjUKvT4sta6B+g8HdYXxmYJ3NLKiZlGdZFm
/DaPe+nv/49gZENVUqWbAuZ8x8JqY6SokTffjwvzmLEFZKLx2fRC1mKClaBeA+gDU8U+rGKgWNVb
0tb9Mlz9Me/nr7olGO8NkCvi4MH0/9BBXAGA+AynOKMp3BFpgLVetCQ6vXXQ0dC+sea8BTC0X0HG
+BABLmoV4WhNBcoRIecJjXBdwy2bvQqM2OfKOoow2meFXhmb1b1N50+fiCcBCzK3a98ytbch8h1j
91T2Y8fwoGBamMj0oFZDQQARft0gzpm7DD1r2vLK20BNfxPdu24W/NAk+Ju5r1ATZeKM50yYoxwQ
72Z54gioEStEz1bQ1vvDmys04xgmKpGCSwT/VXEQfVjJ8TfbI/CmNcDFUlQvCU95HxWvJ9ezAlgk
md6QYZaxzz7quXBK76pM/nEJFjd2pRnwSMx48Rs2JBwJzJsMelCkN/jShKJlETGJVHb3FI38SgPq
cDrP2PoOZg0QeAiPVMK6iuB44VbxBIwfon5+W5aChOEAd4/CQRaHTW0K7Qlya+KXXUIIeJFGewuR
i0OhgozDD+TeTQLAciKvb+NOosHOt9HCh4aQvUZy4CMj6a1ahyv7dSxIT0PEzzbLmSKSAEaKwUjo
6gA8b5d81DgZEld9FIemLPPzGVXYAvVKNWl1fZU3YSyhXEgRvjK5GrCpLIUyiUqZAVi6TUuVtQ5z
NzcA1+akCvVcvvhRpHZPzH2duOOEXYypJbd2Dr5N2/vojernrLe+uRLqGqI2qsSaeaoNPUVfyMss
/J0eS7VbQyO4uDtOoCbpl3HkhycWgLjV3co6w6OJUdw40L/yNbUapjcGc2kp5lgtuagzibOiiPga
JBG4g2XckoFTy+6MCnt3BkPzykTOAXwvrMvza//OPt9Za6/XQwsUIPdl+1sAmke9GdmFLiqxi7BK
C95QUSd9pfLJhOE/rt/sKZRkiTDcPBWcbQNtAqfJj/+nx0xKz0xNf2d4i/MGG3J0YmUFAe3KdYfw
kI1KpgM1QEkN7Hd/5NMbTYuKv1jmBZTNK7PVBpn484rGx65scGVVyAVlMpzrbzCuLpwNOI77zaOg
9Mf/NrsqRwY2ERq4qLvqmDKv66RUpdPz47GfHhkS+el/phVVdPOmWwHRrQZU66UZ01B0PcMWWu93
9MPuNWKfh0llU9pvSR8un8czLRR4liqnpsfC/HxhGqwdjvtDoSUMzG8w69ESec58SkxerJg/dpdC
MoNnMpDVJi0aE/D2D8+ElMhuYam0upngsDVII2ovlIsmrZBLuu66X5OBzPfC6cEKM04fbpR3TxZA
OU8Zi3y47AAaGI0ysuofyCcNtFUlgz3ZeXBZPHjN9vL2cvNkfq1WFwwgf7ts+NYOqaYdN2WfDOsk
/+r4Lr5gjzHuY60GPg2w9p3MgiI4VCQ6jDOBqQ2WvimlwgSTAsY5aBsMn4U10hnrAaWvUAV60iNl
FUmvlVLIo4DD0s9OOVnsRBJGRqg4FgATtpSzj6Q/YiClsE2eKLhdkgRjK2RKMsucYX8XsjFHTA/j
iGRIAqDGPq06eaq5DoW4y/QpO9MCWD3xUm4aRRRw91BGpiK7S9SwoosNYYApIu8N2xGzpvr+ES+u
cpPqBmPCoOJ15M3uLresBL/4lK3IPWWRJPIuG+ubvuwPd2dHy6ZVbQlHAKzRuj2dtiifFWXoKnxM
1s+mbrP7xylzQ/5wEW6rSggn8njGBfVkp5MS8cqin8yTKUauJU5etr92ox6Ke/iAZuCT4zaUCMS8
l9I7Ez+4q9SXeMaXgx9ixPJMsRsqsWoBFAulyO3/beYfaWuUroUpQBRK+n+G0lR2Bax9gdrPsvzL
UuG6QHojJBFbLBIzHC6M8CbFoYAFlAUcQ7XOshyPcR/x7MtTQyU7/r5bEh4X3TflW1O6tD5gD6RH
L+SVz9YBmlzJYK5T//N5vYQCl5YMymI0UQX6pkKKubaQgLzA+7FZD2meERY6O2jxcP35p2Qj0ASz
b2BFViRslbJRBUhG6DyLLqmCMTrkYRkHMMhotmvdy9c83bScPCb3lbdeFoC7c2ou5FSmbaXvatwp
r68Rr9DkJyjjop2mZLLkXGXaZrR4n/35b3s8UQwsT1/zubCVV3QRIi42n7osNmHVkKNUThxSMyYH
BuSCfhwTHE2mlSiPS31tu2lVev/HS4VID+FCwhBTwRDk//9Ob4a8M0W9bGk6FXND4H5id6mlAhiW
HVN0p4TDy+9AuCU73dc/dN0iVi132wGu+7F9OVtxtqQH+2NXpx5NuM4YI6pn7zL8rn7Sk9psLenl
Fn1A+V6khRq0d77P/RO9pXAPb5dj+o9583Y7So/UcCib6TRjT9k4AK2spO9uKwSvgLWPKDHjLuVb
ty86tLD39u+Z5fIzPRkuYaUc9GvjhYqIKs6oWUMXSD+LNx4/BtKBDW7bx5yPoc1IfovzJSMOQoIQ
sPb5+orczd/bof7GgWMY1/Q04TC4sCQQ83goDUEPZdTL+wYDT/Wo+aqfc9v9UcFSdHYy7m3XPXPp
wIbCsDVVQP+gAPYZEgTUeC65YoogeI+6EjqjgEEnaNqYISpceMQSHSKj78MQO3V+wSavFhPVhUkD
e6fm+5oCyvQpIfu4g4qanme+bTNe7TGnLmVX22mBMJ5fcQeqA7vGH8VQqROxGkdorRKKnCLv1dIK
t/mBiZJqM4FrRt8dRMVcEXLxi0iUiExJtAhWzBLHg5zS4fr6Hb0sP/CqDO5zLUtzfxypg8bgzWg/
7rxKGSzedu73NN5E2YE/FbE4+TmsXliquYJgDpH+SWW7yBMI7ecbe1h+C6Y87WzFHlp9b+vhajmd
VohQg32a8fsBDwe0eTXUt7IRBc5kk1V+Mwf6j1pc1YNJ5VDCmo3IgtwIdQUuCMGRHUMyLTuf7u2o
eAkGQ/dma4vxJ8nTGA9gRrbPrC7svmofFZHQlwIQRmB8ChipFleVS7hKizAtQhmuhuSSI9t1wyxJ
Q2ItJUAXnLiNzbYNgNKc5uNyiCQjzelO/1npRFZyyb/LkBlL9x5alX1aHEtzSEznL6T+7ykNU+7M
HWfmZxlEac3e/zXxpRRBLqq4kxJivG43REN40UM5mRPoHkcv60eg+zyf01/yHdt8IafssZKSZycb
ZZo8Tx/F2tMIh0cPsXuK1h6ybT0OgraOwMo6+k2UcKYgsEHkeDp+DDK932Qd8SRGzu0sn0ed0Wt2
2ZZpij2fR57phU/xTup5RY3WQbipDusFdYQfruQrceVqCSEqyDZcM+DXtCQWPeBayrNoEWIOSxcM
cP75Fr/T96UJdhIrzS1+lju5oEZjsHA4h0YCrWHlM3iTZ+XFOlaZbN90SWK2+Pq7A9SjzqyrQ5S0
lDIElQCsTbVz/RopIguPjNBF4brNX3nnYD8YKmOsrkQbDD9GsAS9hskKoF5KJmwEAyvJe91Nv1+F
x2tiMw3keV6WTIEjArqOi/Jt4Hsd9EQ5t0OJpptoXrsEegOONbdDYJJoI3aOIWXsHJpmO9fwKTyD
VWmAARfVaPXqftCGnNXT2oh5Zjs9UkHAZRCKA/TU7Vo3WZNg/xphy6aMHszNmQL0nm1J92Gn4sy8
pyDus5B9uhOUMyz3FjqCzNCG5+g9klrX064prMhXHHmWPU7HhRPvqDaSXXmGOuCKVG3WEvF8dNZb
GIiEGqORVSLVt1UztyPkc3lFDcGySBNWwz/Wvf+ItZTFv3sdCqaXgd2oaq33SiVaf8E0oaxupSMt
8bfvF7ZGoz5MwPcmRFl7pH81Lh/rsJ3MpEX8ykNqS3wZ8kkV6m9yl5OyXVhvu3MZqLOleAGPG/ay
wOTRlYvuPa1trEPaxE+WtEdyM0RpaIoPHDKk1efZlLET3yzZaAjhVkf44+NBH71jTGL1gAgBRVH1
Y1+kIwf1C2CyqBc2FOaJRdRufQUGdezoKXxXD9c0NcsX53c8obmf4V2LOIvH0BEs2MXQK+h0T0Q0
wVKudBrRbw9979+Y5HRx+iIW9S5+gUaxAAxVBgt7yoGyfh3vXHJmB0hdHpbxXyMLohJ6B9Z++78U
hJWpQyb1OCyc3yV1ZA5YmlmiSeNAhGUgp84u1Oe3sVvNAHNEcp7f/dvj9ZgLxsoDN7RY20ChtL+3
tQf9YKoi/s1fcRCB7926yFFhqVsVX8KPJhSx7G7elKC/gxlP8ZWmFXGRXPV+ROZ0SacZ4/MkZuX4
ubRB49qzXuHt5UcGA3qk5/hEHX+RTPEeTPVBdGxZkgPVgJqhfyyjO4QvMXsNCfB60aakb9+vjDGk
6J05riGr91mzTNYv9g317EdVaDbmzPfZEf8iIluSsJ1zQ+N7/jmJLUbQNn3mLs0yL0uLxE+PW4DZ
bV4uRblAYDSjC/fRyRCaGJcsJclZH1BeVFvamAQ3frUCYLJBLL7Ca3XS/WsFTmq/tv2otiiZWsiM
Exf6iH0Ju1BY9W0u4gpFpqtvohzWN4XxZJp0ypeGjcjLAPq/lnjrIvIXXFs7p3EixA6klsorVqL8
zrWoX2YvMNQVdqapIssQ7rtAn31IfwDp08fRlYgtkMJKByJdYd3VT6ykl/472aYh3vZZf4ZdmZxZ
9qPn+qkENFraSPINbu+78jK6Lblg7AQov7C4r3BIyCSA/XP2T9Tn1EgeovMlZsiDoA0LfEaPoo/0
ixnplGCUm+AbPjo53bqWbQpIrfSYgNNRuGkL1ogAGU3Ay1h+Bq+pm9d0N4+koWtBfF+nDMbBbqMT
hCMj39/Bw1nESoIVE6OHBstvx6x2PjCqWrSQ2oBpBqSfg850JX5EEOPYvVMLaYpgHZDYu7Ad0W2m
DNNZKy3AIpunnWomZAxyOeI81af+B+ios6IAPQpik27tTtP5E9zMiDRHeq+9U0T0BMhpHeso8x/N
B7mE5h6eRIFHePss9ctqP+bMma0R4RUo1PFKkg0kHYB+iWjmnX6OUtWsKuV474Pe+7vb7eh7gtde
SqRq9DW95ytldHCGiLeCRcsMCncBZRm66q0xAk6OTdhylwnzynLQGSGajOkllmMx6ofWV1ykHSyy
cgY23P3U35M34RyORqaWWY5c/p1nOOweRqF5O56Jgw68fvp3J2MSi6++JQBnlx+bB06SdSZKGu0q
hdhHtxc/cPW+aGni8a88MPxy+/OKzqF/2eFgoMxn0+I/j+UAvf4OuCB3fItIN0n4p0nxTKDwRMQ4
+4REZDxqjtvX4rix95AWxbVKuBi2TVx8qc7NXAHTQXViByJIBDW/8uNZA40qNDGbWHaYKa2JHRZb
xJcDyp4klR/m99ZfCxX7c1lijo6vAUA9cxwTNg6ny8pA6SMytOS8+Ew+w+l2zNYeXByz0UC5DTkO
P7gjxNwqlM6I94rrk/KMo8WDn8OhatDO1v9VN221Iyao9T/HKO9X7W3wxhgIOWJrI1/VadNpREta
3LgmHK/AMLHZSRy5hQHB7Z3Ofjds6+nuqG3oiB45Y9YbqfmL6sD4VtVaVIFgmsuug2s1YcReVGYw
76zA3SCiLTenj3w/CYC58GsrflDYGSQQkYKE+14t6xV1jaP8tMrK3nPs9qqrlSe5Mu5Pu53fbgRc
twgDhum25+K1c+XN+ksX/bucYJ00cAJHCcpT0+fETsXFGoyqxEnGy4+Tj4GCx0vSXBOB7CQT9zwY
rzuhdcNIvaP+n/52/TBxE4fro5ru521ay69Tepz0+wHjUimIVo7hEUUzKs7fNVmqXIeaRGKR8okS
SWFpwfZLTjMs38vNlodCdOzgNn+Yd3pfAVIWCLLPfYfnB/y5o0jWLBkn1cbsrfcG0R7U9LexvXHw
AsGUuZo269+sV8+zzJpai4fZuCdDaueVnoS0745RgJV5EgH1MPMe2HLxvp1BARgy6GnegRxDUrMX
sDLGicNbDns28nuKWE++Z2rlbsnL6D0POB4MxFZoDmYMC7uomsD1RVBeAep1QbTMPADHFw8lye6u
P12PMbFSG2Rv7eaChFNidlGUFMNaL9jRxtfFbx6yo0l0hfCOmZrsqiAe+5CIbx5u8w0ufLpXkHkP
1Iz8T2AejNU5xXoxrKPmBcE00aOvUNiXGeiovNo4IyWvIHusvpklDvGi3Cz6LxjHwQHXLt189rYF
C3fTSnAT5E4EaqnhuAK+JSAFSecs88vmV9GbYteZNtnbqFgKoWsYJMf5CVZTNTwQZmMLxsWRVLLE
HgZBV3bAmnduukZrEzeNY/2iYReVZO6FbY774IOuvC29kBj8itT/hWkYO5zFZkNmKISxSDHT6x3H
UMXM/eyT6YpoUtHmV9A4XYYOZfdCfjl6IJ/360imyszKjjD2Ko77V0HrEMQuUsv3lUumGOcfX0YP
/+qKZ9p9KiClfZI5o7DAakqZaTEM3oK4POlTP9brj87S2Yo4i9q0w9h9QDABG3S2MFWQqIfWID49
7Wke59rD1IzeId4XIzUNBmCVxXH7sU6jPEQcwYQc0iZXem1X7oeHcff/TtTSa/h/sjV/eXmj/IGJ
mSXMNmqapWuND2goScKhmp2hNOWDIJyc3eZ75DYkIfKg1HOgFNWjhG6MorDAoWT8tzzScQ0g5IFj
qYFH4PSe5XPl1zXt0N2pAVzhl3MhGgRxQCXc9DRtv/yU0iDgLsgS/vtWr1vg3gv6SpeAQHxcv/WZ
PwLclxwTrpax5i42ceX/jKBXRNhQmgbL3Ynwdh0tXArFaYoq1RysYqvOdlBd16HOUmxOMI8j7Xxs
S+J+ou40AeAMijNSnyqhVwVVlOW93KSde04X/Fx/L35GunKNDLJqSDNuOUuNJmZUdERfiGJuEmiZ
drB2ZriRkZkuuvZuEziVtpH9uGSC9ly1MHFqpYlYCtBaunoZ5gCqZQYRJgxSQHCeOaOW7mSOF8Uo
HKnZBnime4Aj/SqtZGwRzYeYKnWlXCIhJq/6fEwL8x7SO3unUkIJbihQwTCWK6qglFi2R6UTUSRh
rOyZdlMK163jaKzHK2td1px/oa+dPDBFgem4+LvMYtrhYYPsyysmgVkecP0DC6GC4H/9B52e3fAu
uyr8v9WJymprP32bJn3+hg11iBbaO/9vXu7snIxnDZJmbZnmQdEvbLeyUDeSXZZypF0YP+28bryS
nzcO1HY3jswh1fRcXqBZaH8DFEbNDX1VNYo+nCzcOEIRVzbSuVLqXnXzS1/rbfJPyeTu5GiywMoo
ceNIeXoaguEvwOywtMP30JZG1YccdjZyAZ4WCp+l4psgANZR6d2oKONLtmU0y2ztKrMUD5YyiUoc
yomn5By5jSzwDQ0kKcx9IZYB338lsL4lVxt2q9tSz63Sbl/dq8ReKJ5f8EByWWoazqI5fKdsLMc9
d6yh6fRxuv4bMf0Y1HDhX4Rc0zIJjHT53SWDw0SoadnwaEcE3ERQ2OstlgEAZUbeLs6rFeRzGE81
ST46WebcpGkR+cQpBZXb2VpQSODl/kxHij/uMfPzPmNCQ+dFOwBYJ3laSh4iporKa2l2WiFyVAfB
FSrCtClwd+bgbZ3CAeD0UEwCk9EVvpNF4vcqe1HdYw2H5kuDKYD1hBPvC8ODKd+moOaWd+NNXYKn
8Ty7IvAOWtaNaZ0+qfLQgekIRQltitiUtk0IzEedG7apugf57AzlItrjwsM3FQ7RnPrxGSzWDNaG
mQ2uyqetUuVWiCtsQWPxOMLjmOTCL0cUtVkZEm0+XdggVbODq+Lg/CHcG43ozQTIw8a3o0n9PpeE
8KW0mz/8iqF4HDSSZpN2Dd5shlqnFqWTt7LVlW5b/j37/CNuryf72V2vbfvlgzBCjUTsyJRE86Hi
Qfp5leJsvkjdZpO3o+O0F7NqA7+6KoJdqi2jFyVznlEsSWiLQBkQW5OhlNC7x+e54XmxleBSS64n
IgKo7IODHKABc+6JOyOPr2/MgcuwOl40yEq9cYY7n+2WNLwGMsynLwT5+tD6uURGXo7BviImlLj6
JOOO3Z4SVJhml/vXduj217mWE97uUw+QeZmdlDP2cC+5KuKwISVkP03NkXvBw1hp/QEekynn7km2
oS1MfW6IjsmGw4EioZS0Ep7Qx7Nzx4ycdW+LxdOhcjz5Sf3JYuICtCBFUG1XTf6ejxpliTkPX+9T
aQfnPA4zfNuSWIJWpbmy6WQGtJof9DByASW6FIFLumqd9n9pzeHvPwQwaT/9AJHAXMTnv4gXiZ5z
pmnagV10fNefUahg9edHhgop6ca9sqkznVexMkoIME+U6Dj6bQgrEVaGbidJTRd/wKTdWTUENEx3
ugFmBjmWsEEMQFgLhxODPSsnB8Y34aywcWthN+Xj0poeXvWRtr67/qp0CJ/IYioaLLdw7i2/B8wY
5WWopDN1AXki5QoBc62+cQkIOI/kyrXKAlB13GY9BSbEhprXmOOY9XWMAAFWCgFTSZw5fTyd7rA5
uhe0V+/peH5V2DPDOHWPcngsscd9V9PJagf3iLRbPGq36GTjgPLNKRZKrpYd5S4gLD0mXRC3lGAK
BIiMVWwK6FQ+JalWfxGi5hFLzFmUbxZoO5kfgV0eUePK/A4jnPDAVk7KgoDNirWPTS21XjwFRL18
V/D3cZr3L70en8clvv00MsfJApzDWyg3KJEo2/By2vVapBd9hKzBAB7f4L5oA24DsuSAoaIVGP+t
8qNZzsbkTxZOJJPBot17qs5ufvtXbLBrq5AqIbC3z5Ft4pOTk07dYy9Hij0HPVjMGgsbA8B49ROk
yHTO5mjCk8BE7t4dD1njGK7y9uSwWRghXmt1t+HUOAq3Ymtwlg9iSNR2Ia80uXrUOrpPvLtNhs8t
aMZjvr8yD9tZR0wA7q3bg/uCbfNyE03KrF1FD+4Vn2d5rxyN9BTqwLlhHYE9enuyeCmfvwK+I8TS
3p3zVyN71dd05dfK8nnemysIu4j6eOufTcwzTwrkZ2cgvWd8LBQs0nx2zaX5YAB0melDYBP1iJWX
wWkt/J2dn+LA4U/nxVZG9ZlZP6PJ+arP72HyXBoa09vebT8TDxfsDWNa+FBQno2Y9zB78ymwa3w5
kK5n93tjob/IaUpoH9T2wERvT54p4cRtya/dMppm1AVIV05e1Q0bTKtRtOqXfRNc9coa5QRMIoel
pIHjC6X6hsKftGcoEvhHPgWTtVgAr1ey4oeRfqZqYWVkDlPWWVsg4nomzhXS0JFHMfPxa9prbzw0
AZ/wkuKir2mbTpCME+42MbXK37lzpz0qNOdTBmLvoJZueVU3tfLm1YD2i6JjNnZRRdQW6edt6tHc
1Z9MwkdfUA6qiMe3XAZ6GHQPgXII/uBZ6O+fsBANodfX6tHrRGuyd/o8qGOCiRGAtp2NAErv/gBs
ZLTRGQjR/i4TOKDSd4k9Pkr62lPzRuZ1lAk2csRt0mMSU4WZVrh2cUp3XrA1HLQ96DjCNCnmN2kV
oX9dFKauoc8el152c0CoPThCAcH2DRgMD2DheS7DHqbZDlqPAb4OjawWbPC4AlZVg3Nqz8JSxjSH
HYyvB+WHpnf8qdIz2LP5nfRW5ROqC4hzyj+KYHT9mVbGJ+ovnsA547uvQHXG8/0rb9UZ+2iDicfY
XJs12HMHUIG9b1AiAdmvugUwdqcNL5YavCw6CpRvqvoIK43fzIcMOgRH5PlAunQ1A5cWXUcfWYY/
PS/13VX0uedFoEoXL34Y394kfrqi+hg1Iufzysw6S8UMKpoMrqopotvDgi0aNppqFPKk6vnBzGDW
S5LgojtvkBlJA0jECSHrTiWvl8Kb5McKH2UV97PVHTzzTQF2Mbf53gU2gYg+daEnEUulYj4HKES8
7WPi4u5AfxR83a8iWv0d6Bpj6oVRcLq4ZxNHWmshclfHnDZAY/yByTm4dHcOVDvn2BVTxYCWSX3l
06mhmjwawOBYry+CMAAhff0JAhH7FblPJB2gArj9RudSCvr3PMR3MUjBw7i9FBgThk4umc6Vd5Mr
Ls0GkXPJOYpZKR7ckCvWhYAV2q6BP20q0F7cDgdVpGjjZj60aXO2yX4GAT8mDdeYHBcKkC+k8/T4
cOR8Di4KK6HWSgo8oSfrYfwvCFdhDaml/xBYl8O7OGvY9aXUupiGd83BU45S1qpRKfB284ZQqvND
DrGLfJWYOxlJ0ongvDMZvhbgaedAgHVLffp9gbj2hc/ODh4ZB7tPR3ZhSNqVpXS15IItld71Suvh
GvEnl6P/gkjS0imCQKvNHNphYfUX5Cjs3c+QAunTfBUN53Aq046OFrxGIx4GT2PpdGSJCgA2kxhq
l4SrcRmYXJ4q3MDmw62F/n6R+siCDd2Hc3jE9i7Ty0hb3xgkwJGSCOAGGZsdgqiVqWzG+D8iW0KV
E8191WueXbGJPJM4WiXNgPUHX9G0fMvhEaxoxeukg7YzGX6dLlh4YFPBXilfpDRF4I1PkHspA/z0
ggfV7+nqfWN3DaEDEYHklX6G2p0efzX6tajOsyCeDPusRg8Y4vh/s/Oog/1cWY+l+iCfMr/fGobd
wujVxjUNRJJyHwcVYsA2op+sE9WXJyLai/B2kN5sQatqjOxpYgaVr9ftDzK5dSah1xjGSUC0vPvE
OoTswGnSuHBvce3i2vlRXKZXWDgqOCVshqjKME7kU6ycIfjxZbAZLtGFVXSPw6Ei3sBSIrZoznlc
QGopq2NFuUd+nIRFjOID3LTATJwcnIQMmPlLnBy1gchdaX9ZgEfv3pWts+OnK1MPR9FP6Y4s3lL0
hfKJCuAJe2eCUiXZbdOkZNPM7k1RVvsbdMnIfCqyIWYkk3bTasWRuXJTatCSI9bjPQW73+uzuC1A
bFdGJtQsSgQTp9e46XMM9hUbo/kuPcW0W1LIWLrKuqp4NOYBoQ0kdm/WPZ7DrOSEhJ99cB7j/F4D
WwCBUM7x2HJ1TBC9iVlJFTYTRrRiuHH7YQXffxj3aqWSfz94Xa83d4SEfysquSG+xLSwIlgJVyQW
cfmFOqtD5qGh43TLL8womzLqS0cQtwcNvntYs/V/Rh0qhPD5UOAN++mu5Et8jyNFbx4DWviDxA+y
PgJZdbsk7Jl4I2dk3DmYmuICIV9K7wjxOgi34r60C0u3SUeo9D2xL9F0IoZRYHMY4eI4fkIL2jVo
+XD6oQ885l6ou4XbbH91Q9CcbmLebByKcciWzvOMIRTcDGu63LSTABBQfnIc8bTBn+fTcFxaJciU
ycjjDB/L40ky2UdyIsS7kW9wYN6RwB4JX7iE+wXwxkLnmNE2BDrlcvNph1xELfqNgtMVd6btkrca
EANcy6e0U/b9poNTSZOtPzj3rJyXv+JHGH/TL4EJ7EsrGJiFF1XqiFu8sXU5SDqXZH7xnkbFhidg
iQ8rjEq7Yv0kiAz3hmfTkM0Hxl72rsebjEXUC1Pvag9assWuhdt1nU6aabcw8EIQUS5Q2bRvsVqs
+CjpirGAZKFpRc8BWG2f8e4levKdwqeYUqcf/Ax0lfyH+J/6ceGevT1VZbbGUJA+6FRXEZ9iicTT
SWcugrHrtVs1lSP3s8rYXfk9Vb2e5onvuefGGQQHTb7RkBAvubQVUn5OqnDPSfSlsJ50gU8PLCdk
pZZuP89gskrqLKlPe3FC5V68B1QWLSRIG/66Jq4sIBu1HT1ELmyMeldnvPuNwgpu378qjyzcuxzI
DQq7IQy96xPX9uFy7KbM7gjftAOhURpI/pHyKUIVLvqLz6iN2HFhNG0NeDVGcY7f8i6gGC2b+OzA
Nc1Js3pn92rOmTOlWtFwP6zDMzgz/ViIbuA5/nayq7AIE33PqMcYOZoGGhZTIoyhzgtnTr36xv+5
zJ1t4a01UcZDsbLJbYHIKMjsQ5U94t2lcU5Aq6e50ZUPpWZHXAQd7YxsvuxLF4adKHiSeBdKwpQw
IJPhdNI5mqEB4GOFRUVLy+FdtDUFI4q8KAHTLslVyeX0eJnrwVMDVB4W5XxpGnUe1ZLOMr9oFbjU
vv4rLSQtLbT1es9x+uRUOAtywpHtI8++uflHXxy84vbTpcK46Ukat6j01G5uI1Y1bP+S2CCgCGIl
fCLloj6GEJQW8+YkRq/JFRQD2lbdWPOgbS2uojOUJRqaBz9LU535Sy8eTOqul3JQ5cPUP/E2QJa8
BLUi8jTY8MP2MrATNUfNQoWP/0mb0wrKio8BcTzUFCv/MturbxHthFc/rh4IY8HZ0bozEGyCWNNm
VvFFUW7a4OTWm0gzDHC0VDod9YGJtydmR6AEKOhy9n4cT897lRiesRwbcSWm1FjeiuBXfVNF6WNa
++IdYjolGV8teZplmSjRRF7+CcS0YhSW9RJl40y4JSEy++y0XBk+bnIrMQVghUfXRHwhkArDazaV
GKAR+T76hpH+XTyxTBmAaWhDMkrtWjsYQi7+Lx5EX1vn+qYtdYXT2H+hCRD959nroFXSTOqM7Cj0
iKKDz7gh7Y6aI6xSbd4YxE+xKhM4FhqwWFW65KMDzcVnIJ1RQwKUKImh/zkv7l1958vTMojaKDDj
v1ZkEEaQ6JuJbkFDEhltfChJeHj5UvSIUMagTPvhpuz5uXaEzLFDpyBNcfO0R2qNDv81iB4i/xTZ
SK8eqMkFLcbkTgY67msAAQAi/lz53LxBVZZhvj+qQlIGuG6jGCTQ6IVmQogRcVnasvfesfulvvw+
xxKmwQakyGZbfbH5dqmz0YSOvw4Ml3/Xf1akbO3/gxXLmNaZxJlInCRDR0qqN3VzuMfaHDBL5Gas
DQSuRdxm5JS6d7UdBPKXO7eKmaEpD+NhL2L7eC45ONhro5hD3TteMwHzTKzQp8U0D9nF+xUir6bc
welA6RhKUi6c+1oZAAgjzT4iOA15PZXuXpMNyYzLBJMS3UUisgW2F5sU98Tw4gMaLae6LFSsZjtz
OSHFrjfBvAylPUtupowtVbNwXlxNZaS32fLzoNrKJ2WFxJV4R5qXbweE3wabptb7yLJoILZ7xX/C
aeEm/Dz5mLNCl+DlD6RRoEPEKSuMdhsBbRVjSOOLt3n7Af86T10ajy+8RYcf683p9PXVZoI1brSW
TarVebP5ACc48ttR5YaPTCSvodP3U1WsjhKq2k69M5LC7OiMaCbmx3X/FPMuqUtWKsXz0498y/RM
J5AoyE51Zo0PdbzZpeXWP4Y87gZL6VwBLGKCVZi7nm+moy5/ZUEqL9ztbEjRTUFlI1PpiE2zt38y
cXNHgdxRUEikXJxzAKtk2oPGCgBQz9SX0CWLrhFrV8Y0etKp81gcoqv6e7P49nI/6O/hHf3Olbj9
3p81+3xP0GTAcPk+cwRwaLvfBBsl22XVVfT9yuVAWYCQMdi/efuXkM2b7Z7xNaqB+Ten5g45wvm7
dHqam75LhTYyIVOBpsbXuKES9EKNvalHlbWugR5i1oI3hYyThPMCobdCW8e3tGfD4eY34P5rUzAz
b9+x4aBYFgS8DiC7xUXCLO4/7IPMpkcimdkrgXsc3wqxPimHpf/jo8fsnZfMl7CRgoXBRTlsxqbZ
1ESqogwBm2rboPNfuKsmziMXiIXJAv3FDJ9rojh48mMICiG77R5LD2f3ACI/z6Y0HNy346jSu1sx
bfyXxga6rhObv5tzNURdgvZoOhc1Zr/jggFn1OsI9MBU7JuK4xU6SK7t3qQRdnvWL9JBFnUIFXtG
6kGKlQtck783uvcCl+XjRVjyBUhbQdzZ+6N+ObP6cZeaMFZYktj1ryVh4v3b90UjI0EoB4TRehXc
HUYmHPKd+AQxs+yHrGLr/MANYcLAkRQw7k2Ulf6nVfVJExK9Fzj6Mr/M+mYQa/g0gXRLAge1I1Jp
92ysU1z7wb/ihYXZyAbMdOdI1C/Qwqw0Q78uSWJxEX5FRRwiPmQXOXpJJNc+9uJE5MEzBgf3WcyY
k/tyjLMjmJYEjX42O3dnghzCH4xC7Zt7U6FdnDJ72jI61SveB3/BBDa1wLSW+c3+YI3pEHoBeGr8
js1MonqpeTaeUfo2CesGmgByvW8+Cm0w+GB79gFl6S51ZyPtfPvIS3Sd+dw+XiZ1TkVZxpmVkrei
39pUVJOWP1hwhSX8ugOlqVqNmjSpbIVnj4VsZhI28JDpIySDEWFUkkDUIQgsJOVoknsqPtWVAAyg
rLpoPue1IEkijHam2TNPtyDf3NYh+eV8l9OFOwsgc69RoY0t0rjDv/GBtZvkOxwKNLulwQ3JcLiU
czulOh3mneH7XYU9I2bK16MdVg5brv7Fetv/kXqK8ohQNZ3Ufi2W9/eohoBMQ82y1qeMpJqHFdeS
njWE4ZeQ5pv3Dm0EaYWzuK4VS2oy11Ll/sj9C42R3bP8rVm6tCQxZWdUcE4GkShwc69EIvZaDPWA
j+fE7z3jRmzMWpqc3grWX+/8WeryzrARTUC8IMZPVHGT7TdIJq2I8ZfDpcujgzoD0vTbhC5YKNZW
O2MG9KgwLKdX/OjAaOQPZxVx60HDkEeOGCSNd49V26MyZbEGA1mxXGyzOcqMklTqN4YaTsiMFue6
WmMtSbfoOntFBMz1oOQt3m4Nl7FKFD7keH8+nTGiovxzMDLV3NcM/KHSZWHwVUDxi+NgGQrkB1It
39xSKJ7oVzwrkzX3vsbKvf4MXsU+wHLtBO2u3k4icLVXF7phrmOYtLnJRsgRQZxFk5TqXA5ACbCX
Axu/GvlC7TK4r5tgAgF1Z3UPcrTpY12noPALtAgnirW3KlGxbUxAZpcsEXKXO9FMSuq+KPeEcF4N
DoExzOOoGbT7BBb+UvE72eKuZ0V29CoPAEWfoviFU2/uOSaXQX16jf/U3WW73jl+MfckKGkZ07fE
t4z+V2alfmR+Slnsa3MfuA+suUMR8ISeHFTgtq/CeZ6cGBaDEou5VmPCPf96hwnUsh1DxnajPCCM
Ji8WXPlDsX2GjjK4uIw3Rf8rveuxUEjTigAu7J5jQP0J4R8PIQrWbhxgk0lTxfATXjm/g6E25AE4
MI6U5AKo2ZOe1zAqKSO1wfc8ar4ZUXxSP0MK2JbxefAzAlsi2uz0XBkDhcJjPRcyPM/WoihvAtiT
QLm6iy4nKVHLaOz84r/kUNS5ypCh/dYRa/58Dq4XHvVsf2qWm0baMA5kCflq0JYr//KsbXVy06Qm
fXRb93K7v9ouwkH54AAx/+zjTzSDeEGT6x3E8TZTUuxsZ7s04lo4GUMyL+VBMyVtrb2l/eOpb+7Q
6PnWAP/Wyk+68KmTP4YNjEnvjd5+7hSxGdGj5+bAzbPaEfgvysWu2xLMYElNi/kR0n/vOQXAALW5
/xAHnPaTlZ/2mnGuAhBlDk/C+VmNewxSMCg9BQQbOJcUJ7pDowQtf2e1H/H+JjikrimaNtdo79Pb
B4WdUgnNJNZUQMe1z7LIfK6UK99n/YheUXvi4lhJ4I39sbq8Xd9ln7LRzEtlvqK2RzPVox9MJLxv
cHSqhyyImOxYjSfNllPdqmt3C9pD68674ktBlvU8DXwZ7GdzaSswJFrAz1OSEjJHoOBguJOsKZVx
FbIGk1rSHLT3BsXIpnOeiPDckaTCs4e8M1T4QeRum4MLZ7xOx72vlK6knbDtQYXA0rz0IMNKyvJb
F61UNk9fxABON0+GqDvtqWcT+rdCtm0oqQsGy5DYP4xwV8Z7rlB8aO6CaVCXl9qinmO9JkyNiWUW
rERRJ84YB25XWb0w6zbMD5PltwqOYz6Gy7NbPiFBHvOHIm2jnCuCoORA2A5LJZj0bcm25c3pucoz
ZwxM11Gc4HrAnQ4FnwXDZUhgOSNCCN9HkkEZRes+5v0kU4Ef8vmwT5oC0j+FRaoWNKUCwsheiq5E
tcISYPoddqFMetUxgscyJABpcfIMFM6tiiMD3lwY9HtqxNrQHbinfEptigir7lRAboSxDXtLmGrL
krm4wQ+mPGf3V58I3rS5oFuHcATjV8k8lP7a5vW70YxAqZ1u6d3uaChpKtQTIFVebs1pLZsyiO0l
ecfPlxnz0s9GzjKOQzVT3qTTEFLCRCys1jsuXriMFutLn8h20bMRCYDDp5NXepc4rCW7/PG6NKZY
AC3xvz3HMriYqiCbpNbOL1S/qpG/Kh36gRbyr5Dvjt48im7Y+T93DGHBrAaMLQvEcglsV8gcxLf/
nVxu3VJuYOXrop/GuGtl411acc5boOTcxVImr7v8F4nVXrtLabyVcyXUcLN0nUI8La25Unl4z8tZ
cjS2WSzFimErBiuOuOw0kHkPaP5yw79GZXVCAPRhXG0jYl9eL8IvubWLBg7VpNFEohFSmwSZGXtL
bDSBq/iMFr1OZIjKZXcsS0D/AjNgRSv1woi32lMl9BOYTMfMWmgX4DYF/NkAaJBbpySYXQNOpGGy
Sq0C/VSVKrlswAwLh/G0RpcsCyRgAHtVDRu4qjW+1xMPvrLEdZIerYB5E/P+vK6FjgUu65GmvdkY
VTNpSVeCJudkdX2yqsDYOlClBWZEwtQIQdwlqfsFrjjo4nkD8dAONc5Lyr5DbDxMGpmltG6pb3Ky
VM+PF4aqmriyBN1MYYFhizyrDOsi5wNr3qXRq0vR5XUNXAb9jKnTOkNAbETAzMhUeIMVZ4RWMKjp
elB+GfbrHW6IGGOGKw/j6thS7ooQ3G8Oav/IkWzUAImXe274Q+oxBlbPcKSvIlc8/0Np0NRwvWSd
2yqWFSgat4AEmS+0TvbwJ1nJmI6VCPWn6A+mnjJz9kk6XU/hl94vNeC23USNuMCUTlnq+6QyO0mF
Q5PWKDCPyK1LGXKV6/vxpsWF7SPxq3XhixZrsxQyoN3ioMRDfoLuJZpLoq7me8XPqsLNTUi2rCjU
7Skuk+PkerddEkvNXKVsmQ5AoKw0hbyZx9bkA411d4EZ2buPjfi0VmmMlbMt8AiFdY6L/gw+WB0G
FovtgheXDYh5bEPUMdy550drxdPiOPJVUthFO5g/+/vAP2gJXnghxHoXIDC6rdC7FBCsBsM8/m9V
EdtCx2vliLfF6NXccQlc/s4NR1DYtrP1oXzmj2Foc5xNAT0JvtCuxbtkFjloZj22XUQnveUujzvB
5RDu4oc00WQeF8HIbaE+Y8/GXWNNsAZbBFOjQ7jOA43awQegRK7WxHePgoHjTvpxqXKHZNq7EYtu
doCJhyqH96ZqsWPaf4PpDCT+UfHLTnKyOY+8X+NvOfUauGzjmXd9DpmXxXOWS7LpClipYxtgo4RU
waVLDl8Zaqdk0pONbp3joLfTvGSVtRHLCTVbHfcRuqjmWTLwDYNC5KeMJ5am1tT4znqcUd3MR43W
2HnMuQYDs3LkdjV1wJ4g2Qi+WRj4ByTz6ZCddQw5njVJNeKT97qT0UmYo/Iu586AIaR74qKE0vHM
C6kN2X/0ZrKPY9WSWn8k+j89QcND0Zz9/EfpDV+ZjddX/l+xphnGkRyh6m+pYzNNSW0LSuCwcvEp
VCsOpKV9O0UitbpBKvkjOaymnJJLgUSGyQzsPTR71wq5GxksBS4QnYFnNX+EzB1viuuaOCO2PvJK
0641hC5AnX1iXt1Dbx+mZzuxNE3GvzeVBIJem5CTml/9jSEjtxDSKdJNaIB6s4Yy1ytYTxJX0pzj
ma1N/cCKjexgpgGbzZQepDxjhbeMQ7drqp/sNfE7rL80vVcOnfff82JPflCuvSR9ZqiAynzURBIj
kn5kyCWS85LH/i9KTlvIc8FJYqFn7H90GHCSaY13Kl9mOHTlRx4xHQQBnYJUXF8Bt7w3rGiwzC/N
58PexfXMt01NhdyFifI60GkBzNIYXZDMz3iRRZiUTv9+N3opkMFsVKTayzJS8PqVSaWUaKZuLrU5
jrqTwn+DcNAs7DjeOP660yGc6rjlGq7aJ8mjKtvf31dlSBpYSlIdal12SosE7+ULEIebZrONSOT3
Y5iVCAazJwu47VyJk7v7A0e02Ud1UgbvS+GGebEU065TMas7AmNhCtHntYp9NPGQp0jKixTzkqQC
zJtVgq3Um+GHK9rbS8WNXfl9pj6jvL1aFP5srHPp5LRrEfv8YLogYd1oPzF1xzPk93DafRk5i36r
BZkhZ6ZnXaYhUbB7ZC1gMVwq1DyB6rsKEAYt6VzbO0koKNSvN+KYD4eH+sahSkvpK8l1q3ZQLAM1
/gk6KmBY1rAOskQLkAmwqWMXFSLNWBmBlX7K2BsJ5Tov+OcuIrWXLA/4BqypChJUCb/2igN4zA6Y
m2eKhokVOMt4LoyapruxEMRTNXn2ec93OCHq4SY/rpQ0a75RwAgLf+Ot/wBPUOquFf6WBoS+hQK4
aLMETZyesuASUy3UNpC7RhhHE+rv7clsyDiV9WzvjsR26UwM89ri0qgzyLflYOqnaZ12nblk3ONB
Pl8/u1Hf+pnd777KD3y0EwlW/4q7dPAXl0qxy9cfyzVajys4DXg6KJVyJ+t7X9kQHW7Ib0zCbDbM
Xi8dDc/a1urqBF8hKmTl+V8+QXdJDccaUXvVIxXhmraCwRz/KArKl+RqphnLCVJDDxRUf6MqADWf
EY1Tp4pSr3TVa1i58uK6GCOYZlg+MTBCjDnTX1ZtfA/eDYfujEu4pRGSVWEnLqg+jbY880Qyn4Do
W7SaetWDOUK/00afQyUJsxmH1zmlsj5pIALoDPXZvBV9Up+7vh3MQ2mccxlVeTwAsBj9RZIYjfeD
NIRSjZ7C36+JGUUMiPo2zcgccnpBnLKnLEbEz8JiWJVZhCFpHuexORM5YmKvxaDaYwleqfyW6rPb
wtywQcYWgcuIEGfYpn7l6apXbpcV6UXq/0YgPHHYAEsedn1whQRb7iggqWyn6lGP3mEmiIpEIdq+
SRzxHE+pe3yOz3O7QZrby7hDSybbI+qH4D4yZUYOuYR6e0iV+y8jHaE2HlsmIwOMAKkSM7QpX7Nd
C6y0/je0j1xMhc6bTlPSnTEP3yj2XzcI5WFhVeuQ0hoxs8gywXJq3NN+mMm0KU9lb7vRayRQ8s2Z
P55aQif6g3YMeluNtmkKgxeO3fJUZbah8MZt1KN4kqZvoOr/NLBPc2TACY2DljrBQqM9gs12ZYUq
OxUAZZsIKVdrGb2XEacaPozl6MgwTxYyc75vW91daCkwE2n0bBXTAepG+AEpd8QBwjO/0A1WPGtZ
nttMKD/rrWeulqwkpn8d4Kbm/glhZCY5Vpo7izGFNZUkMrfn3D6J2vzx/l7Grv92H3fqPJnYj6wU
ltMtSRgj6OXk0n/mf3PGsR7Npzt3xXouZEKd0wyqN+VxR0u7MobpkWV3/GVdP6QvE2Iz9vPVZ/yu
ZvhObh4mCjqHLghMS4tU7cQRVLjAg/f+RXkaA5iKj3jgCeW/c94ihb7qVlqgTYLVNA4qklMrTY5t
6feIM5GejlndNbgh1RG720dYCVGa1tV7EJ2sWyxWxQnOHCSWAbEQgRlJmLWSv2x9KriumgicyWdU
nUpaTnYs2tzGLMUMwJZFRnXQ7e9w+vLf0x/lkKWuO8kpz8LyVSp2Y/EjZWsiGGuzUUu37GKyFAHr
WQT1XGirqiTBRgMg8KbPdrLa4y0EHgAxITjmvJBnpGyfwn4IeMDR/rlhuxlkKaQ3DmRqvqvXO5ck
qXnx+N4qCXHY+I2kmzdIBByRdFhmK3+9Bd9NhdQD/fP8c4/vHEYidgnH1Lejql63fN9P+UAjJDsp
+2LTqV968sllOxYzB8asC+iVjzOSH2LGNk43VSXe66cC0TRSNedhjbaK+Zi7nc/Ld9wMmHcUrzpD
Cw4qHTM71m20VTLZnQKX7iJ4QEGWgfaANHUHJBxNgUZrUDY6XlzJDi221ry1/EOTuebaMKMMy8tf
KbOAI1B+9jlLgws6hjxoHhs9HViVkN2ejik8Obn2xWdkLbPSLlA4esm4j7r1rpPKm0KfxPkrKSDP
+l0Ue3UwTq84DepSPcFjjJW5ZZdWps1TwoDLGHVfuZArR20JDCrNnZY++ogKQBnSUKO/xaANGdfN
S+XDojHtQiv9leLp2TXahwOC8qVxLcWtxtSsmyWLu6AVfaY5SLspgdUfAL4yRpS5ckmil9r+ZZik
Ryj3Ka2P448Nqm5R5lOORcKQ60HM54q2G2efq51TsjzS09lxtM1Pni88eHZWKicr2cIuG0g/vbSq
iGWZYBAZI+HW6Py/CFnTVLKMSQdosqeAZ1opPxB9dEgPbh5QiQLCBadFjNnRHRy5E+/sxurdcEQs
VXSrsG4qxT1zHDwVctQ526DHqRp9nVknMRNue5yCVk20FWIybHPAMWRc9Bmi6E1E+d/dfUMAWKIH
ORfVjhsuKkP0H0QZZ5/mFsCaVAx9Y83Z5N+6pIw2Xx3sLJ/AzsVRg3wBOaUvd0Zn1TMXEh3j1iSr
7epV70w6VXf58eINhVWKt0fXBfHNFu6qYDqg4oA7WvGH3QHPWnmi3++XKf8fAJwsU8tIYCqWccHV
3jkDobb1uLilOrzCoEUeVDPUsZPe9qbJrLM9IfwkBgj8eX8EM1j9szL5bYH+wvL29HuWrBKbAZvu
/75nE33FM//LuMxJo+BWchlBp2CX+9tZWhxdkuP6B32zjAQGg+TX72Y1f63zoz3mpx+FBYMMa9L4
EZo5siU7TYmCCPQ3PB7SBCjOkBFJhPOp8Jpz0xrnyj/+fQfC2ERoDr3sAjLrFj5kSPSG4CzLQaGF
pAysPijtc1Fp5meDWfHkyaXTPMvRNgAFLBZOm57K/+Ocszuhiixusld0xrbOXUQpOgxDrGmoggxz
qCLtpWnVeb1qagL+Jd5kuDX47FKDn4vuxXPaM0PmaFO3t7YuoAO4RX30fRPB1wqi3XXd3gpWAZlJ
VAXUh9QpWS9JF/pMCHJQnsYJ1V55adVdDMN2fnkKUoLnC6P8LxVHwevF8WU5h8rixbpGuVmDVFZc
c0EuyUvi2NWDHOElo24HAueQ3gQV/U+2joRwqbTiEVmbzMfYRAkbT6c96bzVIsoKZHikOT7IR+dQ
aEubSP+NsFAQUZaGy2U8EJARuXztySp/l3+UI4kNUpV9O2B54y7qrxKPZp4LehRqgRN3E87w4WxE
o6+z5C+uuoGUHKH0k0ipdJ0u5f1WMd72qeA8xPB/J+iuQ2wYOtx0MLP5rM3d86MHM6HiYhBnCT+E
Utyt8IUZwEYFbtgDRpXv/fsLo5Vp5NaDkiK8US6hMyjXyy+JNQ0CW2w571uv343FwUJuB/J+Yizz
mr8tnMiYyVt4XJtezJiWW8qUKF0qWJTvvjq/i8JsHtZ8mc/P8friFYpQN1j/SZLeAQ0izX/gJCXB
q7D+U6oXz7HK1yk4qZFawhc8wWnt0UBsYzIoAvuB4iJyt0J/U6ItnJtzT9xaifwDjwA+wD8TTqeG
kyMizeONjvE9ddoJeRXi6rv8fBs5oJ0d6CkM7pWRn0EpnNOCiNkoBMJz9psZPA2+/s71Z5K8v5ww
tEbUbFzdpV8xMx8TwZXzklNEFHmmkPOG4/w0TmVr9+xWEM+kQ0LprE8CJU12lVn2v5H9nYj5KTuN
+WR3aLg6PdVVFN3LjVqFObvH2Uc6dnrp/EVOKenzUWyWRteCSWrEgbmuz+Bc3J5gZr2Bmt2pe4ul
XNUyCXFVdaAQ3LYq6k+Ah5pDAPpg3WSIKtRZkojHQyUHVkvxjCG8WALNktHwtn3r+5LUwizdNi+t
GpB7JEV9E+iFAIVQszcIb+xzUvTvEB0tuAfPoTYDTNf4cIEausaiOCTZlANkd3R7z9Zjozm0bS4o
ou1qGoOfSIZ9wdAASeV9eupInIlcgi2h61jLiCMHtX+rioX26Jhiq6ZIgyj+iVnj9K9UgcA0YWgt
wWqE6pIfypQ/dvwc7bp34gD6yawADO9rfMNLHtPF9WFn1IA3TnVvKcnfY5kAx0kQx/Xsgi50MalF
Nu8HtdYhjimc3ENG0Lnmc3jOSKizWIVDIMJgL0WjAkU38akGPJU/bo1uwhkE7LCZuy8dRxeybP7c
1oZjAwB3OpIu/nhvG8urtOtikJy7T3c/XmGpDwsU7bdo8z6r8KAtHForuMuTmfO+4Wr82ENz14c9
KUFZUZdFCXUINURMfilgSjiUWc4qF8hkZ1TAEftm/OkTsJlJ5wAe5Z4nCHFmahD5b0dbQDlrnF5M
DECK9Txmvi3rmZwr9K2zBk+APMEYr/AN7ZZAtIC5wxf+zcpnprRw4glmZbTn1yorlpUtPDwyEbeZ
JP+VkoBgRR+SHdrwvFJJ99HZXLzmmda/sxdoO4WKrYh+5MQ3nKMCCrtv7NgjFnfBXS8d3s/TEWn+
p6xfmJWCLPgJct7IBtWnW/nC3kLsl7s64NEqYulFk9ys7BdxpknKxUowKaAD9bsEn6joqNQ7blcx
icxllXFH1t5VlMhGWYnaVQxx62HmLffOMEB+k+Rol8+d7U4jE0taXSpD422T1a44gVISHV9f4Y/l
lNRzmPucqPuz79EXOU32Mfo46a7gyQZD37mPkOn+8w8V7HqUUDAlanJFF8NneOC15wtXGEpmKTue
Atlb6XRAopg1UQrsZgdP91QLNUiprtJ0lHHaLcsFVHVXFS3cteqGvOswQIvauJMd3rzRLOwI87Ac
/FjPqvskk/E4FmTjw9Mp9h8CVb96dE339zz4z4OROzjURR6cYlPR01lVOc8lfzwd18AVDAQB8VNm
AztFGHJxolqeEEhlp6guYDnbyY+6ogkLTrv35Ixjh1qKAOLCNoApJYbrLHYMQdMw1RBasXPF3Djv
kzJ8fvUE+5B25IdxlieJ5lKG0fItq5ma7D62KjJMGxW+4kNQ4iKwddJm914kRaO7YVQm10NeH3Wu
yV+NXGTy7R3kEU1/m6uvzVn2EmU069eU3ta3ByfwvFxCF1jcFR7yC4NBhDTdZTuGK2y7svSkDGa5
qHi/bI6YfrbAtgt16IGVpC59GPS9D1YoAfDiTlB/KM+u2/7lATx2LSDyIpNOd1CSg2SzLopIDlSc
LVDjdweR/GjYojV/EuyBk6SsoUuFFYt5q8wySH10PQKVfiGQ40Bf16feTuQRVwnDZsmPcePf481U
AMiM/L4r0BvX6dMIXwRcUklK6fXP9Zxr7SFQj1cf0tQIc6TAQxX2WHd7ib9LPJz6/DIgYXzobvLg
UQE3KlEnFCyPtFXb11DaRmkfgFtlM2JYU3x4Jes4hPPjQkzqhhQm5BI9qu+QVEBH+T+kW1vpYWnl
AnwLhGgJL4qcDzHNW5Vuoub5nzFOp31WT8+2ZNevlJp5SvRItyIJJRsyjJuzc8IorFKwQ3ITbav5
LbwDfd2jI4mqnf/mXe/45EVd7rB9OvYrtONffkRCXmuUzbwYktfbOdbcATAIHA4viq4/QB21FAhS
CHX5SC2Yd6ShAVEF/5vxxajbDKTb1zcfbeZxm44YRopgo3/03ILG/q+o+nkLctRYaNb950ZN+KUA
ygG1JaoSr5Ejya7DMnrzOBmPfdc000hAT7JRSyBOl84IZgUWm/D73c6MFn4WZUd9RczVRwEj+bGn
Inxh9t18oqaMClS8cQCEh9BwSv7LdyJ+XRV3g4c357bjD6+zyYQv09o9yG/+puc7fjIwPVEK9kI2
Hi/F7sMQCQYwndL5JasSytxtq+JRYSsK3Oa4DHhyyjR5ery7wdlwq8tb7bFxOUd6WVwipHrKOCVp
QWOJD1wgOdWDMQHjBDYeIYv4QvUMUZuIqf+NX/7nH1rR6bR1FdxCXLEt22ndEmknyi7TE+qqxg6P
lqtZqGkTX70QehkOYdcpYXKkAb0WivkFJknfAmabjG7IDvNXe6Utfpx8ZxeZvzraXdzHFUkZpveS
BMaYgXdgpPoggQR/saukgvGnAGpFawn0U1EAl8N+1icGuF1A5bYhc7M2mz3rF0XVU82RDjkc67Eg
fjOP8oeiCsvKDjc2CoI8m/oUqCsgNSraCs7LSFuWH9jBmBlEGWZ4fxMup8DvCmk0A1kLD7iUB0bp
kieVvHrWnMk6MQsZcrhYQfKnBSaJb/X8ApzL4kmRrum4dz1Pn57WwJTMrHc82+WDkvuaGxADVnKc
+sMM97ObNE/cddCX3Xu0JyNBmE7V8ZMMDgjpApa7sDR/szToC5K9oxKLHxEFU0cvcP1JqSshmywQ
m3rs5aeXeZs0vZD6A7QP2Y/8LmAOomUse/N6xb1wxz36TJgOGYkyD3hNVnAtjBP0HEONHVB0Kmpq
f3gs5UBnsenbSTmRnRTHsbdbPs3HDPxE32kzO6xusSY2qvAdRiF11zGHPxvbyvd0mgO8XuhyAPCW
UhKj+Hf4+9htzXcG/TO6PSYkk3+DiWOdKMlxVZv+JFShyggLgME5gvMhx0fkxnvaiT2frKVHRE2H
UU+nhCVZllSpvZXJ0ghCUqBMwD3njWiYML6dm6b/l4D+3G1SPjw086gaRQc0YVZ1C12mzSXkrWJY
15ywz/DzQHdy6ERq5gyp4eNudYUm1XbA/wPARkM0sYhQYELfBiBYh0/p7TwKwMOC37jCt1QcKEI2
GqxnqLkB2mmjQaawTKknBxchNiml2XLfiT7RfS58yqFmUFxsbRii9seM0N3NxHFHVzk1BV7vvg0U
wNw80rOjQ9E7fiUbp8pY/slZdLhzbr3fpdKbphzHpIEHvJ/aE8h4K+0q3OnJqyWEfsQIOzEd9OjE
014DP1i3kBBh84bV01bPJJwSjIvnXIIol1qETUxJoQ81jVAUvqaBGj/tYU6zuzDvuHectSRjk3y5
wBRysY93E+GFETZEJoHLJLtUt38vL7toq+WvyX090XxrOEcIsXgWerDPeoaMLCU75xi2/LYuEAyF
wYEupH+8Blu+TxD2jfS1mSaHnq8p/d01gufuPXMXvMKIt58tdaPfl5/Y19nK8bf1/GCoaAsmI6Sq
MmN50QWfc+Ekd1WKIH2BXXDNjkGeCs5gewpv4+h9TfFEbTVY5EQ6yei39stlax1wwpvhwg2evBZo
Kp7CLaUujYEsxux3BdbcXLNB471c3sMiHfRCqgKzKXTh3o6goAvcFpC14WsPNtqa+gVuWjH67NUr
SDUdbjwOvAluy1jj4wcVbNqRJIyneJ6cHQ1xWVIpDDwrOb3cX4WE/CZioE4AZCZLCWXQATQxR5uy
9+i/GLcytUkweqBLso/XIkvLDsZLc6LkE26z+Ay5hzHex6d4sHlFnew1I9uZqpJYBNukYw/ifSDq
gwVGP8Eom0e0/Ie04RO0qkTq5yfEii2yN+sD/aRYXv1xqSLoEipqPuXiU3yrA2o92B3/1s5OTzov
CZg2ePKk6+czpsGBV7oMQfBWEnriOyHQlW9UHRFZv+yjlwcPU0IYFby3z/J2tgDkjcKanT/QW9lc
yP7jaONksJa/g7UuBTxbV0kfE2Eaa4EKTJueCy8vF70oV2Urfm9Alk07E9m1BvFVlyq3iVmcB6PF
bcf9z25rbKyCdXXNN5QJJu15fPiwSqXiH4CNce8Z+E9wYHjIfohLdzcyhEDmsUQlc0vd7JyyGiLU
NHlD1iwANnvwNmvwcqruaizcp8NKqMiw7G7PmsQ5BSOgo06b0B2BAgH3hGy4+ZtjH9nRAcp6P7hg
cL5BJnGLd8ZAoKaKfU8vVYDJKPBqjxGu+2K7F50tsF7NshgRzAumYaniQsQk1Eh1Lbqc9VxrriNv
JE6TZML9P5lAp8qOQ8XZJTzMDAb4fKZ2OD14rgSi3IdxRM2bV2dDTEB1ecc4iuHXn8sL3F4iPAEr
FFAYHRRnRn4pSC2YDZnxH8HHAz8VQ80XL2DdpGx6N8/cbkQcrvPiwweShuHjV/xUHhsf3xxQ9FfK
AOMMTzqItuPNnAxmpoOOvVErvAvEMyLXFhtz45f1Gsgxe6vsHdTgzujZcLj6UBgErQUBfLKcGMwk
3Hw5D1Cafa3W5Ls4R2JfjJDMXKNnQNA9sg834vUAvqDBDNZWflURwhglwYOGJRgvEpdLQI4qfRDm
qMusnECbz739kIdmBiNMNFjqbYFDNGdzos8OxnwjwuJ71cSwfet4TmTpxFJSaY5+aG8MqHyszwV8
eDOlQEiYej3/V1KNgv5dxNOP9GuwN4E75dOyqW2i6JNdaLHiYY9tPlBDCIFm+SBKJ8rfSmGF4n5l
nMwi6kk7Gj2iEBGm2IxjDvYTGIt5AED8TwQKj0I0h+0igJHhF25jXdjVAszOZMQYZ9bcNrQclnhL
dn+KZa8+itgJZly29NZKjAx1bEoPHYx5+VX5Twk2Q1LpCQ1qlCJB2c3fdqLqJ183MEtAe6iIJFET
efDFpsxheLK47yarHxfztgIkoCaIF/TP/LV9PxbnDVyOjAL0SnURKnhbZT4Q8FHfN2BwMvC9HDm3
qUuk2GPCKcKWzr/dYsi9YKlEt3+RYsRCwIBP5YnhBFwPGVb5XxSgLftrwuAIGSt+LBsgON1w9Yo+
5JH8zPj7xeyz8oJ+WgiOrxvLhafcuqsVXG+iorsmgIvrMNyfY1LUy1aYD5pcwNMtua6x5iF7Sg5a
PX2qXbmIPw5rv/9GnUMeZZmBsTw6hI9JrgmfnKLkk2Z2ltR3wg8q8suLKXwmUAt0+qnI0AE/jQ0Q
KSan3ft4BRh95Dx96fRfE8lnpLsLFXqa4960l+PZDYvWREYZetIrpPhv3beoE99CfbDtj2ig9njL
11EPdXhwhkAGrG7s4KxoOZnjwR9XAbFnpoff8k9QMWQPK0ML74aYrsst5UcZIVAfXcMH9xGiBLPF
E75Y9xKxW7wsp1RgaEKIW7B16YC7IIg838JqeJPxzSPIPU+XMIjY/drpF74GVVwlAEXphgirEF7q
XubzmBzH9IfXROAGwDIzZCtzX3tkaxWU5+oEIJdva0NtemzMvwn7dstlTlw5z11P5NxFoBZzGzuy
dj3j4cE45IDHcm5zsgj0dd9YU8Xlcdi2zy5WRfttiH/NvM0CEiRPA/ky5YV43fSqPsZGi6m2nsT9
Sb/tI0vALfc4XvyMVZnzpGM82JJ/jlUXpQbZcvoocYezIugXM/PgSOPPvhutaK9XsxVWkkgEiXwp
cHYY7ujiHvd5jAtw0+LS7mP8hDRvcEGU0PKUD1bIyh43NxOdq+yaW3Gbahxxy8OM64C0GdTq0mW9
2xakaGCNxVCpVhRFaNZj1wNafA5R5upvF6XxGIn7NgXh2O1lV/AQfuMRfa+hZEioirdpb5sUcZLz
0cs37chhbOlTwfmPhdYBtmsF1RkCKOWJLqaiAL/XuKUMB05gJPPy+qq8I40jFAoKT81RoH2Hh571
8XVmU8DGIjD2Rc8lZ7WuxqZwoL9xUqBmIN4LfBKboEC5LoEkAI0OLqdWup2ihroJlnJQ9DWtdV6A
yKP5XEIg7DU3htLirDVnGrXnu/ABfr9B+CsJZLhktIl9r8AVNbDDX2FoN7kAg3xcqBwF+FGdhDRH
3hwpclbqcdFc9OVm/bDEo/39tHwCEpR4A/pZMYyjZDPwcwHLyJibGEjJnsYrjQSeHjDjVf+CNQ/Z
b4bKFkT0o9DyqAc+u872oFshxMLfe9sc8AHA9iUBy+vqVaoYJhQxQqWOKcWN2gcXVvU/mJu47cDe
8LIp9sRycuZDRjV/uwEMboMA7phdIQcQdaZKP/D2GN1vHe/dGXEUpdedxshgywWB9Lyy/CMJ4tqc
UBGG/DAtUG/hV9gAjIOiEK0z8MFG0XhM63lt9eYwPP37rVsUeSw9/k+xhEoCv0h+zomZ8x68MakQ
uIWytz3TytRenZYnvAzA476DmlziDEgYPsHH5VCvEa+Haov7VMr4rg9/k+7EckDuybnbnmkeL6oe
sxGJKEgZos9kdlZQbedSLFl5/iFdurtFzHL9CMIW/wlI5ZUmcnkI2+w30GuNFtWK9rGPeeBd/MQY
+L2tg/iBSHUExGK+wIWGzz4nNR5jpCzpHOeB1a6RdxoobcXkynSW4JVZMxrjXY3FP14OksNm7TXx
/X2EwzYFTXSDcPe1z75JGw7om1OSuOOg56pNCQENMLJQ5IaJqnkS6I6AMTzYrsR17K07mkHopUyl
Cl3oLVgZPGzu9DmL6L863StxFf8poiPlWGpKEiI657tmZWOvEw1Pz5bzVFqtHJUrEzl2mQfbCHay
PiVSkiJjc6lLO4XWds3xyDe1tS6Di1USf+99beFK63feJnjXJTU/401a2TPhcu9p+P2jMrlbqObp
ccjN0VLgBlLjAbGW/aSDqf/BUsMWmcbGCqjISE8RJBlx/bV9yc3GIdJdyreDSIl/v/VQbvmS3xmr
DTbvwNkYwk+ZJQwc80crf6I0t6kNCDzLyNAmcunERmR+wlTX7jOAkVFRS7f/7TeoCsxNuoyk9vvS
lbaPy3eb9uty1OHVDcjTvfjiNx6gM1+x4A+Yan2tyKujmQzJ87k2nyQlfdgpDGyxQIjoxSAYELVr
zSHkdIjI01VDolYza7+xVrsF7CDbbS51qbg0+WzIcnK5LUeOoyKbeI+sn1NLcNzh40+Iw9eJ3TKs
ch/8o5uU3Kv0sr17d/qTe/ZhrnSnQQtlRFWfBCVFwb2AhxheFran5G2jM2nU15ccVgBdSQaZd570
l653leLMv2czPcgL3rKfBqF3Wvas2VYf5Yt6x9D+sCxRDBDdF35tcbcJeSAD0n+OWArrHHN/QA4P
HfhbXsh40AO98vqE340gsRbyiaHGLuNr5mCRN3aIDxKl4WrlckmVu86nm8aAA+tEHQzAD7xk85qF
u02td0xxQlBKwfCCLpb7/2vfOHHRfgg0Z+UFhu+EvdK34Wr5Uzzs0Gn6qhVzgQgtJ8YIOUeLbeEN
Jk1Af8pSYlNKwB9qWS8n9ktYLLdw2yAGHq/XtSLzXoMLmhzELmqz8oYZpFcpbjTtCDGJuX6syax8
ZW36/NZo+cCVyHdZLGkd7HOErRKCCaoR97iVIIdN+mtlobHyDYUuz+WWLo5s/M2WalMuTUfnLV04
UbwvoT0OelWCRhmZ9/gb00ek2dHYV9roMX8TpFga8xraPlrpSQA6nTZ2hSe4Mv3It58+c+vtTztU
DCTrx1zKKHKqh5mn0nlnj0m/heM3N7ya0xq3Wk6BNEllI7VNTw7XfzExzt4jSo8BskDLlE+VvmK2
3TJec1UBrPY6ZV6Ya80MaZYoS7C4lN1dmGj7ujZOUaz+N6kGBD7d1AKmIsJh9Crpl5bWl4Iy8+Jm
l6tZXx/Uzx9zrgry73m0qhinmKccF9UC89e3Qtvr8lsJB51yQoyqAj10kgwVzIBHyiWVOsK2eDpn
nJ8tAwBIn1DUb0G9Z7Hf976jb6qw7U4PuAC46M6jNIZrKtNiswNPjvc/+IldAKfGpYKGLh+oBwg8
O6kT3r8AuI/6j4gwbUZpr7jWWPFnuF1CEga2iVaRnyOStK1YuPdxGyoPHN3Kuc+TcxL8lcROLErs
4o0baj0Hn7fJ1hL8t2+1P5H+yKLyqsQAJRBfTtENa8p+cdlYqcBnCcP+cv5s3mXzIteRCVwNwmpX
XNgLrEbT2kg2Eq2xpJhz7KGoVLht+UgpKtb1HqXoRv9g1b0MZhyW/h20qeFAMjzzax4vf5Jfee7D
2MP/IfJT94z48xLWPu8pmcj5leIM5Yb+hyY4fIq/BHBlMZ5HVdcJsDnUGv5UBoj4uqx3TabLhbzB
9N6jg9CcNfUWgqO5XS7JZ6yCCUvcIWSY2rCVPA30eMD+haU1iXDlBpTA/X2M7XwyNZtCsslHF/5/
MjwZhpd+GMk8SKqXtL54WJKxc39CU/RAn3nZxZa1Yz40keAXOQBxuAmZtKbbD55vhRxgDgXWQT6U
9XjAbEjtN9n8H30lQ5W+gZcESc28f7FTO337jNP9O7BlcKnN4ofbLIuPxPsVa4mUE6Wf0gqZ9gld
mYwKkEMCw6lf58fJ3JEwz5ttVuqkzU7cSkaI04h9LiPL3QcDSWcnJaWch/ZrFwgema/t81bP22dp
qXNCUdFZEl477PizKx6ePpmTcATltV7rKId9w5YB2Np0ilVpV2yEkpJfq78oDVS/S3gKQvyx81/J
m4G8gHLBguzI+p7zuSmNkExOHYe0BXY/0ZQw146WVHQjRlXRBdYPAvMyQfo+J1q0TzfCd5U5U/K4
VEf8r2SuGZBl6WNRToVl1x12fGt7iErp7b4CObOiawIlsibkMwUwy7OSFC0fIGZSIs1uZq3I2dzT
8i2bEfflakJQt5e02yFys8G+C6pEZ3mnkLDRRt5ey13Wf4yIfGApvRBs45ralAtHneuxMtsuhjHK
p20CGkKHUEOcfdyEITeYR2FgGnuo/vOzkGAbK5+S8XQR0ohmDuThGCTBHzyeJOnzmOnDZdb2BpsF
n31BOQYtr2LetqcxD+c9jeSLPXl427oTARSUUrTKbU5GNmLdf1UFatiD+rp8qpUBpJ8FCS9V/BDh
8Z9Ac0eriEJfB6tg8CvzPniq2UiIV/nv0TaL60NElHr1CiIfq5jNiLICmHQaoZg0fSpqvZQzwtq+
CdpkuZ17FCj17etjXFcQoru+MynDClO4qgbHiVa4KIpOesCEscnimdx70enNkioNxyt1ffabB42U
KQp90r9CSb0Gz2hyi80EAmB3LHpsbblbkHWqWAk50nxiy+SK5F7DTXrrcVGqitea5wWLT1yaTayw
wqDtC/IVjKj7F60PSE0MqMe2jIlS6R7TZYJhXOIskAGRl8fjWmLNQXi3fb4pf1BMZShYk7KUp5L5
NopKQcXRE2OJL97rYbcNRad8tMXSFttggo3b3LLFTz8xGtUZwRBA2u3C+tpmWUlBS3kPG4Bdk6qW
ySBOOuuL2dIFoR+tWtOWBYGb9ikGwMtilmAQcePEzTfWuee03QybsoJ4dtyAAItzoosmw08IUP+u
QqP8MTBKhht9KRR32oJfQQOo8loLmWDW5MgBRLSkHdzDv6jL9B/vPlr3XP21tTDSJWXYrySNz+bs
SWZtmVJYpGno0nhEpfCylpVEGNlX5QXUYG1znWXwN/EUWdBgc6oH8aY+OSUyFIJA5+KDDIDjUV91
GdXByV/xlfQ2e+gt+IztOIC+myhUbmJbJynGqqz7BrcYiFRESJ2u2DWf4orpPdvew0/z6TU8UWt8
ToG8SlyrZrbIQ4t7sx9aMCXGjeVP8XJAYqBDdwTeRnApWsiJpAEGAO36DctFPiTkkG/uJLlGjZZy
usb0N0fmWLsVaB3WNcmJGZ7PuHJH0Np15eCkf7le7lzlU94ohBrj2iBzeaIEDt2unSHpb21I77Pe
8UPMhw8pN8c8qjgIDt35jjGDOOv+CzoPp3yJU1yXrEoTGKOPyQ4aB2rxXu87wByY2eYp8tUj2SVC
oAQrzUTAjEQp9uFyw8IXMV21uaVoioNxdEBg/zBD879zrCuLgmGqMGc4y5xmTa/iOyQmMdKD22kz
YaRm5jTxuDIMaQyZxENMwbKucLpvVjWX93/DsVfRYjbByi5gliYVEThfu830nBauj5bAeebbYnp4
Jo/fon9XsOJst42ZOSz6+m7pv7NpQ2cu3n7yTCc9MYH/WCfIgd33ARs/lH7mzgkCGvruhkl/uPgt
7uDn7oK/eQv7UcZ4nuDFntH6DLcz2j17dbGevamy6Oagg6cWqCmVj0LGBIocwX41If9L/ofaifFb
V6iN5Ykmw8EmV2xwUkILSy0bco8ohEFyOti0eSqF7PTv+fGE57USG3nm+zpQkxUlntinjTpM/6ZP
4dLj2a/bYBPJBpyCD7CPYZy84bILSP3kxBQ4l0o3ar4b+knfd0j4Z0kMUbVtyijpB/3U0AUcM215
R+7exU88dKIzaFxBpaocC0cSA/9z7wn9M2DlloB6KdFtQauSLtWLbPUrj23Hf9gZ8cVy+WSAC07e
lX6kH5I7fAvMw9ARfiDpONPhQZdoQ9eLLE6PItzrcHdPfHdU2WChBJu7MTXipPdGm4UvVrMHYL8X
IDzKEzy2N/4cz1AVSWY5AcKJhSADDB5gBPbMLP1sj0lbrFrf/+xyiH0wme3eS4Wsz2rae/I7Tuxb
k+HdlXRB1F4RRq70aLRkUWWCSstwrZFzlZf7iCvtH96D/2O0wkqJ8WbG/CHW+cFvMdAUxfhNMZib
8MzZQyENuEOH97ufBMiFkp5/ePP6r9WZ5LoDHGzD8LbQpg9UP5NneE9h0LfDIPkBJy9gSKBvLv70
81WdykULgBi4fqIYKiSzmhAbwUnmXqhD9oN+5FUFt/Cy0Oxi6x1yLuyNPEVBp0GvOvPYUw1L5ysJ
TvtVa4dt2y+1DUArZ9scXvaYb09kSKxPnLdNZQYlZSzkxPuDCSqtfISvv2pkMQkDaRizKaP7hE/z
4jI1PwAqxd2YJn9YCRIc129MGlE11ODcf0XSR7Pw8/jLkYbPb6uILecMOOA2RXN2Xm1FScfukDPA
sm89oeQRKwp4FxDWBJx5I86Qd7OD2043MYfLGCCKuGXp4F2jXs6CJSE/zFZSZ6CC0IluaaxiOL3Y
NH548S/3w1TsK7hlan2dA5xQaorfH2Kff1aIhbby594fhi+PCUhGE/vlMgt6OsizSHcvpzwnYrBG
wtJsRDUjMj/PeGXvSnMuff+nrqtkf16ZdYcMA0LfEBcac3JcP/0RJ+n+Vw0nXwMfOs74yDFRzYqR
hKCkpJakh/ESkDZgOPiEc9Q+wrIvtXqPFCP9tBDy+6NOTdygfrUuFFxElmBQ2QU6XWqfNmwT5rGt
yPOzPoCdNRHli2noWY23br70x7JA2GL5DynsC0XcZWVY4GWMOHOiiCNGVVQ3toBc32A6UqkmLNn5
3CR0eStdD7zBCqvu7p35ukbP5sAwRKOZlSpi0eaBbjqdXTrtqxxsTvuXBdsFa0Zx10D+k+mvpnhf
2FIRa2mStf3N1V+02QssMZVAGKWP5RLf8upHOhdLZvNBNSEnrJBtvGQwJhL/LkaDnoNvh6iBD1Q7
dlyI681U6yhcWoH8DjjYdz76X5UoqHHqaDPbfRCzzRq4HUkcLGLa+9H/4Q6qGWs7tnBAFo88JnPr
knQnJtkS5bMaxXf3UaXQEEvYcJOy/yxyEPdQy91uofJM1I3UGzze86YwYorhjrREQVQK33Ahumct
zLjG8Zl+xvu6F7Y0DrUDuxoqW2VA7hEihxFLomEWqEgLNXZ9RZOt2A+Kd8paBrDgXuHLRs4rNLE5
HdpaL5cNjRl+FtRSfb36za7WvvhkenHR4ealX4lIQgguCBx5tWW26xWvRdRnWxcdjhKBL4jsQ3AH
bG9eZLCO5gUYa20cBvPSDcZiXmzBnZwqz3GAcL4Mnl/qXA3zq9KpfS4q8CBhKa7Xr8jpR3F3TfW+
ms8yBvjRgciE0YrOFx3/RctYPCzfXBES+LWgP3WJf3Dt9TWg1YKeWT8Ksry9rZDXSWcX6z8FqmLg
8DH1Amy/vWDDtQ+UtzluoZWgigLTO1J5Y3ntMe8EU8yEXVvILFutBoRAu7GDczBHBb4Gpv9HbeFW
rdQXz6+ehOqX1WXt8CnPffUg2hATiUpFD2y+QzLkvscY/uA08bi5h4c6lS+K6M9n80UL9jOiDJhR
+AXxgKjf9FEOvqC6EBazM11TMgtx/EXeOXhyZzISf2eDSeoVzpKZQK+9M29yXoNKAm1+TATG0TfV
2apbnejVSAKnn8Ia4mx3zmTmwiEdCEbvTYm6nPSGmrhKUlngiVeYv1gwtVxkXpPWFFrzw4fK7rab
gVxjUd5A8KwWZPFAkt7cLCvZWBLdjRbrF63rc3Jl47gihYM1pE0cNDfQ52jMsepyy1YFn5P0IiV/
VYxqnDdtXAc75o9hI961rJ5JGTdnyETJRQpWUmoaMYjhmDQDxMxyA8LB6W5jy3Hwhi7DU0tWC9nQ
30i9N6dEoTBDAGKA4/D5ZPdsPQ4AOLk4+gcaNuSEh2Us/GJhMq3JwiicGDklT65IztyKeKnFZdkJ
CbuiRbodiXB2oRi8r+8V33Qedcl8iWfZOIDmAcJ87eBnnxAWbNq1rvQJJVX7BznleKoeqyoooN6r
VMZ3wHgKYhYIKrVIItO76RHTPdrpaUqnJqID/zYX0ttUD22o6QOW2KM1kmyApIxqyLpbN+PHH8Mc
paD2z6dFFStVVgtqnUowFYX+pQ4VY2W3IcYe3bGh01zKyM0xsLetiJW7KQYhTgoYLShavIpR0ltK
EXbauyEsijZtv0zGhjvNrqOLWvcwMDO9gGRnaxMdkxZaIQsUiHdL2cWoy9stgMkMGh2YIzvGfuDL
tRCc9TSmT1YnxaX/DFll5+twtnvyj/qr9dIcwvLWBE7A3JhHJWNbfnpM1QqkfdrxcxpcUgH+SDi2
RP3zElA9MgYtzk2/vqJHyI5prcqyPqIDgr+KEhYvIM9H2LW8emVJePMlo/8rz+CJcgCWSbhRzj7A
oA1Oy1cI20RO1IJyot2anJ24rXJlhTYm9lCb05s4OcOaME1xmssbE7AuyTkI2IJsF6XPEisBZfHF
YdvXzTHJrdWQpwOfskd7qWHSYPdF2Id1Q4dPH8CiAnoV8EDx2j8jC3t7I1kwyvsihyEo2eOb3Jte
ELA9Sq0hgIimkmvhKCpUEDhSS38tUOzVnZOnPv1NzTNtSycoLFKTyZ20ftWP/uCjIyn7E8uVqn47
gOMLZZaixnMDX3A/k1O6Oz+RdqTTwWKI0tBcLqhDVq5IdqUGLOiDVMtVMZXfw5P39FVtoV8KFI69
uBhhAapy1WIVhK9G8LTGrdVCXnz6z5mZ/ahoVb6kZZqeXRRR/XUkpOAiLMWbBDWivJrRwZtBncjn
vhC6d+ks7hYAZzrE9mdnFgJBKHP8rMvVGjgbhgfkGFsSsPxUgdYLP3jzoIRrVot2lmHl71cdRtYw
VJ8/7MzlEY1XqVVApZAvDxeEd02j8AmdH+vQStrwlZxmzfwoHva4Z7kuBT+LDubo9QnMoulCABCW
kWF3mU4zw2MxN9AA/GjCD+G+lBfe5NhPBkRYUFL3ETW3c1CAJwOIKypeX+/eULbVsZZQkMOUFrkG
SiWiLuFxpEW+H1bgNyoHMr4mVr+G77t475z5ERJiN6iB+2VUUirowTNQViiqPEwWUuUCD0Cqunv4
dGWgCWyF6Lujqa3c1gev81HsoE6VID9uIwwUDzIIjJBvmm0iCnRUMLVN6N+EqmBy3TfY5z5Njt4z
vnvTUOKT1/9Qs+KgcxdL7s/cIp5DGFc735qP6CNzMckhCwWYId7tiFZfyl1kqVLhVtnctn8YGWi7
tiv29EMYRUGZTwsPiBYrPaAdZUJid+dtL3gp/AcO3V05lLihn04V5KlCBiE9fsUkiirFafEefKJ4
QM2wRjkpX92mtV8+yN6RqqcG97TFCYa9kARTziz1iNGOyvh/TVGnxwJukjD65xpBERWqfGCS4Eyi
B/DA4QvdCGRgwqm1IHG8qn/TGm4UP730bp73VzwEd8yldX2BO9KU+Mv2VukYAxyBBX1rqcgHhq7a
5I+NbKa6gIcfQseqrVKQK4ZtduoquB3I83tSoaLtRm6HrPwFjHouvRoVePHZjhWKK5KQgDTenGkZ
HU9wIkeN7wb3KTghGQHu5kVsN8y+qvoxmIlDAiV0b1DIL/QP4ADM+/NPy7CngNcBvxuClTJlg8Fi
28vXqSXQRAxvl1CclVZxHfYoZL63dXNeoibFWT/jL9Tx3jwxgrd0Sfb8oUidDxO2tTqbJuj6q83N
Cd+YXGEKEek4Kfp89tL1jz1Z+DBVjMU0Y59iuNo4ufUUcv69s7orrCgC95+IRIpkFm6n206QKa5m
2kZdi/67b1hCj5lnrw8Ex+lg8jvielPSruXjyy9tXh2weR+22FbWrApFx+kVi2dlsWuGNrvbuUb8
PtuIXCMbK4648Zd7dFbNyimmCAE/RNe6vjBTMSM/41V1b7Bo25oEYmVXf3SiKHlAgnq24EUEpckU
8yq/MLTZ2aL0A5CS/JsWGl23BAPGgvd+tzqW2GSiNTicE0abdOAsKb/umD5gajqtH3Kw9Jty1WTm
xNQl9rBwf0EvVsZRd4+5pP5x7Rh7HLb8PQlzv7McQO9vDmBDId1H/xS0ZSUboT7MR1RrcqqH+7KI
/xiHUc+AhZi7asCJzSF2ECNrvd+6PO/Vgg3K7DFPzM+WyYVY1IzEydwbA6QCKUrJ3iWFbUKkt/uH
HbIlrLyaOnuq2CGQO7LGd+aK0i9s1Aiqiq/eZOVNKfWJVa1w4VGWNjiUYQKjJZplbGcxOGlIttZw
1e700Ig4OMwNGFphtM1ItgJP40+8pAUJmYOokhBWNCZeuDKb4VwhaZ+h7sjJa1EEp2n21PHX9iP2
MQZHooVGBWoBLVvFfPBliyONzmVFHJYH54vEJP+V3Mza+qqBRoNA8jo0qejeqSc/lgvumI2BoPKd
dqUJ+8X/W4LUaYEfwGEIH2mG57ovPtkrwmN9NnywuMiK1/EChBpIqQUG9eN3f5P1ojIkmgKRJtop
T27IulMknxS7m7F0XgQRVgZQulxcd3JxhqznQbj1H0lJOPay9buS3YxKbGVELOzIa0tk1r+Wns6l
SPROe2j/Dn5bmZgBwBIYhngEgF1Z/Fa6KatEnzAQaF84ykPdzP7zKH4QgIjoZO9NC0KaWh2z6U6w
1jMWcxzxgFsfvKTEh9/EZ/rWH9zL/er5cB257RFr60KVeK2FBjngms10bdo7j9aW8y+mmfmu/ZaU
WhrYqBWZunG7Ty9FSOTKZy46Mq4GsCnCfuK8SLnjW+VqKmLvrmmkLglzVdo+oEed1Z9V74qHWQkx
4Wkk06nUd1LqA3pIa3c5ZCT4HohJpG3vhxWx2G2Hay712YIOFh8YiGZsjczzCAZY0yufQY8x/7pL
DaPejBCIVXkOflslxaxnu9hDbMgdxNGBuwhGxjERBn4l+fHdYhlQM6HVpKopS1uPDVxIsE0WvTcP
FJAEvT1SB+9m0KdsysqgXr6G2hhq0Vz7mn3wRQ//lUjotpii+pTdkYzaF6wRecWCILREKLvzd5xT
DcLovS0sLix2egrO7p36te3W0cuFZv88nN2ufLZGtNQEt2gbEdS9oKt5A6VOAFZ5XlD8CphIPFP7
zMha/JovTaWZao5RTyn3Mp10rtbfCbpfeGPB5s9JyW9fNJG8P/N9le02kWM00xmGxuOSpvSh9GH5
e67tcxc8RxndYdYO1ulQUujIud+/1Zaq1i3c0vzdG/6ODgl/gq6zHSlaFVguMZghwilqgiJj6zMT
Q4bdPpXIGsTcPGR7pEO1LC8UKHvqqewJ9r6uXT8V60qwKfmuPXy/LmUZkbW5oIy8/0/Q70wlL9H1
5IxdqUj1EY4ZdAYI4A4NHNb5jNZbfJBHgfTefNzj/XM1P/sPIyIBhldojO83h41as7SGttL4ldBc
q3m77v4iSOQrrLbPDwgCIJwmbpVcQNLKmyXBSLaZaunkxISZ5QUU9bstfMfHocnSATatJsxleVc8
CuMJf+MtUiKX1WTja1Nk31MJh0IqLvE/ngq5F1Mwmfp/BtGO4B1fkLk3aM08ZMhMMUHo32k6Ytxq
GgFR+gEkRx32B6F9P4Ty2loOtTy5lks3Srwo+WO4e1ukOnNx+CvZnHUGPHTCSY2F4wqxRmhd7P74
R/NeJoyMK4NHaBVeVTarAKSieB6+BoNV0v00Zz5DiVRx5rxF7YIL9TzqWK5KSUErK4biTRc56KWD
K7A74fEkKpeWvi4Krs0smr2P5jeXy4/vtG+edV+HR02l4UWkeAyxX+XIE9uahyBUwmHOPi0+0jlS
kNgaF7kjMbaL4m8hcfW/VT9yEGHEdaudzx0BGnSuJeM/blOB/yRTitKiFm0uHnVFoZXuj2b+Nnpr
QLf53NLIxLop1jvcmOQG2IdNYBrXAsofkNar+aZ3kkF1wUFbasckq5STdDLARKFkecas1KSobAOF
tv8pRYo7QBC5KyNX48ARungf6Xuq1h5t1S9MMFp4qs4ONG+2mbayy+vdNgR5pbTEsSCUkttwpyeC
PZFJGIDI3fY4F0xLhclzkppfl9UPhWjIAyEIVi+DYXeJUS8K4eD9UfvyZJLgltGXe2k1iF+AGitx
mXrsx/lPtHkfj+4ElEALjTi/ZoOnKmVjb8MuCFdjZLAdbGd1j60HFNeUzusodJyMLYW3AJ3pUN4V
V9pZjEBnYqlj9k04qdRcSbocZglvZAywxK58fb0RVBjPA5pVJzjXNCJCxjV1Y1tRlY1LSJWwIHAb
a+EQcX+VMfIILJQhah6GW1/ItGNFUewnovbOKMonY57c/w1fmBefzlNlM6xFc14AmJt8wcW3FKQf
LkLsxBxJniIsY+Tm39X4mPQ7EQ/ZVVp6zpgsMUeG0IU23kGn+kG4zpYVg28E8DHWfwYClQlVKezY
O0n4NKyYwIVjCOxKMv4VzdXfDei0sYD3baUkCNDfqAd8GK7bj9hxi03SrcUu1jgppq/5wLFKClqs
+W9KDVKaSEwQYmjPfQR4HJKbUE1qvEgVqkjnn1L6wrX/kEBP7QG4R15EwrvMz2Rfh08efiiWk5pF
ifJuLPxwT1mzqBO5Mpd6v7YtrBhqBIX1mlA6PQ/6btmEMwvQNa/0wP961JQv3xQCTNMnu0WDZkN9
99Wj8Z32TpyNKqA3b28Y6Zbzt8Fb5UxjQbi5eqi1ieGhqclHwt5InWqJaQd9ojGHiqmEnAVowm22
Qqpa7et+80nCjiMBdxDF/1muflHjVoIKz9N4YlQg/DLSi5XSq/JnbcSOdpZqeP+0zig9fE8THcIK
JWv7sWQm0MwMx6NtGaVSEWL6ugpRScrZ8WPLTwWdLmUcIyWHhsravMJDTQ1dh8HL8nqKbqCcMgks
G+wOWeHcQMw6KNdiNq6N4ZtceweP1bgycaCr8AxIVrxSM4/eDEbjUo/n1pGVygm+jnZUOI9XvjdK
9FMctFXb3Cp8rzP4Xe3GD/hfuSWHVqV/Hc2hoMynTnBA61UoxYrehT8UfswnHRurOZsRrp0HW4Xk
R2DpTL2lxYNomEaccLLgNx3FE1iU+GZmprAVKYO99G9ipK5UZ34Axz+isgidGx8crbsdLDv92uTP
wxhLEz50cEi0D2eYoNDXk7gw6+aHEA0SFcLZ1TY7GR1LlHgYiwU5HHNkdq0ksiX0FT11/nyNIvq6
GcJKqp7x68uN7WNndzUZq1aAP9cFob+SMazgLFxZ4SJpwW7O3eHzHsZXf6IBx3fGC8XIxMwninc4
rnlOUas9egPYI3TZHjeYKD5FpR9EC6SkQTEgm0+0dALsSUQilfc/0Uish9oGYTrpcLsQj4YZqQ1b
/rlv3mBwjPI6gVvjO04bsfunu1xGlaufM3aZtcTcX0OOoup9vNxDyoNdpb9xoCuPOqKS5x2i0d90
HTPw3d6Lgo2k72Q+764tQuHRjKgP8fYZIZP1JRy+hfsEhZ71B+QayrbHchChhWXkct853LelgyJO
Fkiy+XhR6VDKiU2AkE48SgfSsEubcCoRt6FUyiToV9P6YDIgO/whgq0JSAz7wTAPvMhNNrYLSyj8
xTDN67oB01apyhjLCxwR6KCE+z/v59tJv5wZk4moy2iaUiMLwvvUtopWE6CwsegoQdilf0yRSXi9
lWIPOvFaJEiqLOKZ5htO9eLd9FhJWolOdxasbm90d/OQ62/E4lTSqX2s0Ng2bHMqavQweIwZALLg
0JrxoFHFzvkD9EYSeCHr3sEtgIn9QHvhv9grKcn48FTp4pf+qbBxGagV5SWhDI/sZqxtIWY5SKHJ
cHenDnAlTtMJVfFW013Gai2jP+H1lK+rmIkies50OnkfhIaUpmNOSt6uMEq0YCfo4biK/DdvMx9H
Ku7okDOO3jUxIkb7VvpSfvoxfBS+JFYt70X6qsfbqhgKqhDfByvrRTtzo7IDdvUjlYWoaXTWPg3m
ExshSg+lVjTVFxTR7Np1kd0GXbsU6Afkty7HuuyXf6tYCeucCC28wAf9eXBu4+etd2JwX+iIlawB
TjV+KkV4t4EphPKULnzuW7WYfun7vKqCJQsUw989nqQjkqK2ayAVTN/nelIPIu/nXrnoXhncGgAB
HViMH2GeXMQ3k+vaXMmPmwHQ3VVIL7Yi9al3TSYHBZ8yqAEsyl8+yV75+qy+sALvSZl+kO3kUjUy
wAs8bRtHnKgGPEE+JZoVS1Ao+D+3ZAS9OTr73Jzhy8G/wmD4GQaUpYWeul8ZwDJ3loLvnhFAiZhA
Vx0svjstyuZ8EZYohRSjgfE0YIBg+b/W8ki/ZM7UkxBh+KoYRoAP9nemH3I+bjJnCUauUIwDt3VT
fDxaCnJ+PBjgqpaxJb3WfVJbGE4Zh/xdlqrrf8pRQiAhSNU8gETdJF0TFLJWrXS4zlS8vJDZ1G7J
QXxarZb0lv1QRhfjsFXgL3SvsCrlklgsJ3R7waDIrBLo+opgSVDRuZEaY4xqAwMb/B6cZ+mK3ZlL
oubcOIhWZrgYNAkjR/oZzbHq6xDu6O7Sx/LBxQPg6ym1l680lZTHNCnl5IZxeXGiNIdsaY6FUG+S
ybpyZLYSEHhNNRguCD3PbK9eXOTmbOYbWcki5o+cTy8nvqgM1xvI9qcFzaWuVriaL6NLJ1uALPfV
GNoI5W9Ty5nF+F76frm3X3yTCSx4Zc9FdqvaeKx2kPeU2s+jYYeplndl3HfFo+4AWJpp0NISozur
CQILCrI8GjVOU9dgT1D5Pa4eRZWrunrE46M8k+KGGjh19EkDilWwMB0e/APD9AJlE9J1bFg23zk3
Uf6Lw2Qg9jHLdpGA9L8tl2cSHmCFmZmqw13BJkJA3ImEO/vVO2RvU1cvE4CzKiLmgs916KWpHLNF
Wg7b3SnHXNtLSVLdWy0c0hrffe3bWqpvSWjOdmXNI1lH7ijBxQ7m1O5+MBO3qx3JG6ihpMwKC9La
IF70ws2Ed1zEqUlYYTL9X8Zf/b+JhEyktUSgYUXGru57UF5Zo3jXxbFnXzul457W9nmr7LuhmuEI
8OyIe4KQBuTf4qZHGhHqQu30yxWvwcgbUvUr1I+Mdkk4po4MiTrBQ3Lm5D22AHNm53+h5eW0B7JZ
ApALizNghMnHpBL3zMdfjI/F0LSlIXS9BYWTacC9VsCle6N2NKCCzjVL4IX0/jlSG0JbdMsyFVRk
BWyA4gnVBTZCy64RCeXHgUSbhCfEjoJIlPE3sG7G4ilX6R/9MYXIRh1cgku07PUPlG4Qv0sWTPw9
tPGrvfOuSPaecEzC70uKKIbBAhB505TcL14g1cvjDmsRpskbECZ7whrrHv5vxfq5kw5mlzd6B85m
XC4fvAFNFVTMDx5z4FiTnBIpaoOJlglTDY9hWf68HagehUMCJDSKWiwlCb2OuGcH97L0wtQ1fD/A
jCxGB20U1YlXY4Gni6UUDSmHqBcgf/VtoJsLk3r/yX5I2hfYboeQESjHg+MZiFtPSmNZERNSXv1L
RHuft84R/4lTtaIE5potu4vFQuD7OSdWcLAtgXPq2ccLfW5RviomqSspCzSkvJctI9kTGL+NF9yw
lveHQS+YLeP0QvcSIxhi8YICJGSqhT7GV31sErsQsQ9x9L03C3e2ijMH/ybtad2ojZmRtBY4H5OY
9l8Pb8hAlCEnia1K8a0MYmvV7Cti8jsP3UUUhVQm0vN7V7YfNCsOhi1Be8DvLIbxHjrQ3gb9XlOV
ZM1fWTLzofmGHipxg28PPXuQh2hE5WwW8YuApKrj3lSX6fRGEBXe9g4k0h2qHU20kog3luqEtlrM
WR7ng97vQ9DC+egze1y8XY1p3nqbmlrJS37EVSWNZr5VVNKveu33u7ZAAX2ZW/3L4PPDw3jrO0Ug
nA80fQMLnZtV/QbxeZ/fy580K5Hm5ND9wY4v/vgLiZnpKuJXp1ysw8UXgb3TEPc4W9eV+wIwuCRm
Es2r7OZ55zwZUwoSrCu6ll4Q4I/yDgVNL97EHLVuC3Btq7V3f6Bz21k5CbhU4yYlPKXZMaiUup5O
XyTgzQAEtjYmmtYlNazfAx0Fdv26cBRXHlEtGMom1nEJn9PhLYqy/22u/Bq15ZCvQ7H7WRA8iQPz
eiG7G7ZX289bFDxnHmHZ3v1RXZrxS3V2CrMB77JMMLM5CQfSBcjp7WVzLv1qXhNSlMAC++A6DQwc
psodRhefAvky/7ZQ+gQbW4ICmkAbg0TFgA9JYqoqh6QF0NLe4wlvijHS0G3H2DRgp/aBYC4AXB2Z
Jb2y5dXhdEh1GFfUykt9NCPwKdKpA1Eo2s0BcYpF0dO7l7xcLnVRtqea8z8jGQjEGTa+ny99uu0a
a23oq4Esf+C6KdArX1GOevaLw06J0PgqsTUC9v/yrL4b2Cxw/VDIiVSvgkFhiPwXGoLBOnkzN+gL
J3TUQj6e05deUGJMZtK2EC/5neTFdt+ztINoh3VAIi3ThkJlC2NCyaN8HAbLEGM1ekevapj4n8Jr
DAqzr4Qb/2y2GGzbB+UVSkcARJaqgr3eR3F/s7HFjNPFkAJK+UtJkQ8UymjXdePyP8OimgflL9eP
3X6LKL7PKpaWWguMvmst0BhZHwrE3M32Xu8vQ2gav/P0SS6O88XMZfknVYKuM4kXxMcti/DA7HOr
diV3SLaEJAdZTXoa/S3RS3BHf5h5Mqk7GVkb4JGZQVFYiyK8N6NnfYXSVQpAi4pcetxSpxmLNut2
F3FvTlDJBSkL1bvGbt+3m3NncCt30Pxf5XXEInvADEuVarfxQToBZrgcnl9dsApgw72h3h1/5w+/
Sguhs/G8Ysb7Qx/xIGrEz+s+rCgdX1/wyamtrCRXAPuBfn47qQZBhxwOUPKzk374IDbrr1ccVDF+
d6t2i0Tz/vFt6WvuIpneq82oChNXyhSbFSwCz9C/o36YdEAOMGFS/W8cNkRASlz5HrelKpfPk1Qv
apEYUx/qTUXMULrdvQRFtMeKAUUHXUJwrIO4Dgu9KoipmOvWDm8pxcQd/rdaJCdt44XzANNa2PlB
EFDMbr+SzqyMz/MuJek5ceDcRBAkmF3/k2WOAECkGi+cLncuT8PTqkn0A5QKziy2OkiCdMgGVD3g
N6dNNWVlPDwqKtMAHC1PExKMrrxsFeGJgA4rAAlKFVaXqR4YlGchRMmaLhf/SzzR/pmR9MW+WGu3
7rH4Lw8JMfPuCzyx10+AnlV+urGDKuLzkKISA6Kvg/J6IeOyG+zzttezrtVcl7wk0sm2Wfky/Vq1
nF6ZxJw3X8PVOWATJCXXUlwfppWxT1ajJ47S3MglsERvu/rMdzD2XejoH0Hf37M++iNhOQ2LrNU7
vrITu8LnIXjVXAa+GYcxrwmxEsPWqPfPhZeemghLLny+l/xBxEwh3iUgfi7MRUQrujFa19rM6zJP
/aRFXxdwzo4WVgKN8s0u3liknIp42PZFDA/aqAQh+Y42DtDpL8yThlab9SnJ7qeW9xwgO1VZpXkU
fh2tL4mOwvF+mYgUijxEfbXFCkNJuj7UgpXAHL30yToaTg+h6oNgt8OIGdLNV87IKLtKO3KSPmh0
NHBsBbT3OC2VfurKQPnbmQA6ZwElTj1MbLpkCjBSgNO8Xl+zJzaCBEYycfltU71AjugNWoTvDHK3
JO/JjXFty2m/wnfyH03YY/LN5uI4UT0YHGergeSokfxJJHnoSN7EcAwz+m8IytC0Y1JlRpX+VSQU
VMN8v+tJTN/oBKOu/fqM65lmp9wnKe9kAKIlmYtSE8mtk+TwEVPfEALjufsZQq4cNDwB+5+6st67
m+tmirju4Amult8LrxkgK/nsT7Ze5HARqbEa/qjK+QaKhTBv4K9QYj1MSAgOrUvzUeTZIsU+7nmE
7XNwiXXpqLldjIOIiyFp+weolynt5GTE+kezNr1bX/lilelHdYmvU418xUdn1U2NI/dH1Hd+6T52
jLTcXX+NC3FkVQmeSkvVwKmazzD0iM6P/a/LhZFOGcVy/FmWHOAoPZdJG+C4xRAeUtkgyITt+oZP
2xmba+a3ZAuE8UpLS5suXkz5h+ufPX3ySpSl1httY5kmAR2AcvdeGHyoQpR0puiz0oVBE4YK+SfW
0DQrxDgPyK/9W59xwLwD7kiTR64bxQEawz/UgzpUFzi4E9Dtxl0cAgAo3xqe2JxKCZzglLtxi9Oj
4kQI+O9cL4eM5Y/+qxY1c7rZ1ddMzA6qJwEdSZ5ZStAaNfWNAfw9MwqEEggMZcIHTDKMIFLo8MQy
c8kGKGbbPepQV4o3fsE5hwvG3jEaXAGQXXQp9S1liB8eRhQaD4DwIckIoiefNMe0Bp7flUkA5VX4
boGzV+87oFhSqZDk4Ag4wII5PWo4P4jppyXEgGUCbkzju3zlYWfzO1x7h4hn0eFbqZBUrz0cBKmE
mtuL8YlK/yoNx+I6LY0VZsMa/0E+qTyKA2qiPtXt7QyNTkA10PN27oU+RX45bR51o+4jiySy3av4
QUViDgIchh0IuzALHH1RT4ovwJDBxClWIj7Dz+nj2A3/Cn+/uOd6m6MwLu1RLLfWbWoio/ZJCO1e
aGy4iW5dhZbUda+G7kjTWhYzEZustLP0s3jO3W6REoqGowISHiILQqnQWy+K3b7sjGNioblxIdQs
E9mN3NwFLnMVSazwUPFn9RbnmhsqnlXUFzb+gyBJ4kC7vO8OW/1oXM4KTUFL0iEZKDJbltiZVxfn
bp4YfIYFki6UUVsbkgBWeRwsTzChbJfmPvVJlNQpiJ2LfsxHZ551tj3Y0MZRiMrL9rddl+es37Wf
+514lltF5lCYlKj+QuyOFUtig9Uuo08krK7xaE4CsmPUMVHaHErz3PCAguyMMi5d8Hihf7cQ/EIT
xMaGOBinBa4LibSVE9uRgQzn1w6Ki9oVKbzwp/F/UFVIx4ql7XbKA5K0w5s16kOjvabIf/kVmNwb
WUl2/keJCMIqu8SDKrKRKuv5K1muWUe0cuY/Oa6PBNZW3bwV7outQzDGYgiEfvdOJ2o+PaYyiiD/
eSPD1DIM6bQXpEhj/77MS8pdw3jKMkAxrmVfrETh1+y0FQFln3MBYpTWccbTczL6ojtStEBVdtuU
FMfUs3vGVEybUWPP1Jfx7mCNJoZQ9Mzp52pp3PAevfe4YZ6o0dMFMPS0LoI4o1LO/g93M7VY5CzF
QfyzY9140zKIgb2oPvAu6w76prDPtKB7CBbVV2g+oJROhWhOXiKpLwY7RjeiGgGyEVbcFEJ3UZlE
biKuqdyC71zRp5mIO3LMxfVCS+Dq6oGzj7YCshlF6tjOSvvW68eBs/xFYWqbdmbSzBsBQeb3Azvb
qVQ4IfiB9+beEgMJ9Jo+W8MTYHDsYqp4zGUSZI0eijFyKCwMAvzuBfTaDgVkthUwfqsBzIv4dJ9Z
OY08Ui3BBz6XlnkGRzy0O2B71jZJbIHxQhkdtnlQk4fnhQgQ1Na0pfuz7B8a6iUesdHgQhoDGQrI
M7iVHf2Ohrx3Up5zDPN5VtsrZgOgvN3Was8iftOD26MsErZ29Bh3W0HtOT+DCgD6O8qlF+Nbe8Xj
NXaTX9adS2GT8LraXhuJxLiZlrqCajT9U7c59oDzsdJlusUpcK6XHBrAsVuueCA67WSbPuN/4n6B
ZCVwf+difVo8eq4y77eMh4iB2CKYJOYwBiyKbiZM6zaLj5ug8gU+9AFyHsSw/aBb34rZJ5HXUxt8
ZbaHJ8xy8XJ0IbN5Fvrdsl3xw/AuA3JBo/w7QBPneY1XHBAq8TpOoSPy7vNk6ad6Mia5u53T9yH0
7z/w4XJMC/VLQDOH1kwOyy8oZi3puKxZVjnGFtotjYjQ4E5K7JtLmv0V05y2zW719oupHKSkd+64
Sbl9oJ/UIq32V3okkg5EtetANSUrCJ8i9fP5+Ybwi+M8250gQaG89wRE0q2qOoBPUFzGevFvxHKA
DDYnfGic62V4nCrd4tLX41wC7EOcx0jXmYg1W/EGjHbe4Cpb4kJSQM4T7kpSpaN/w0uvOM7zb1+Z
B8qhdkuRZtsN+dvFYFOBXpFiWmzIz2800lh0m/WWo6Phcx/EgjlOqIAhCk7TGJqqJQ+UAY42U9BF
ce4tAvSCWwUJ4fMhR/1uTeHw7PorcPJlTjvIUkDxUeVK5eHK2WuFpa/7hHD9utpPuP8ocX86gcDl
4AfNoIpW2Ppq1Q7aRXbk5zkYSrnTR28dnfHIJN8lJ1YXiXOFkvMoe7214e5Q6HMoEeMvghh+h/UL
JFOLKovcN48Uu8EYMIXyWAn/qYExiE0zSWZ5ylSHD2aoTSvboempZkG7JAwbKWoQceITPzwhBGAh
VZGfmAi5Lbr6t29JvvxFEVOQgQuoFyF948CM35KzRkM06qWunnsyTfzJzjbjR7GZmTWTLATPTftF
JKN5lkMYK0ct4RvuXhPipMOJ3CLIESjclp+JjWfbyK8VwFAq/PxKrkTUwS+Z1OG2nEefzo+ijaC0
6XbD0hYWjGU2smV1MRfvMtUpxztCsdKDxpIHmrsDhs3c/1tLgZb4G5v76VU+m60P0V7QDlM119j9
K3uHgtQ5IIb6yNv6vMKbGhtdEXg/pUa+KJtPdEienunkPy/u/fIVaevt05eg9t/Gj084VAob7ZB1
JJJveJ15sG2eNlu/5piXBbXiYNQI8xtMrNqOL+Jix7s/AuWfA1+R66tX4M0Qle6OMkq9N2fn25Ne
trlK/cBKdlbPlPAsIDHGkL60XsOoOcDWudXKWQg+1lSIF9mkGasM9qcplS2pFXY8fQCm95/TbZLy
RF/bDPXXi3NNIRTWXkjK0BTnGsoYK/4jbif1SChmzzfpV5rQl+CYnOjsld4u/feQ915SGqbjH2jn
Nu8RrFE0lEZfQExErVzbGdrJHR4wMyj35xfZKFm8GYwiuvF9ffgy8rPh+rUpLYy41Er/4lec3s45
XHpJtT2wvaXUfZcyZy9f0wPIVGb4PePW5krlZ4LceswFcxwsAyfmzfQfteX9iL3ZnkbZ5NCmRFrB
DmYeNZwf3P/kStoW0xeVm9ms5AktpFc8GdvNIeaA3BBi+XoqLU/2K8Q3spml6/+u972uK2tygWmy
E4W/zzao0QHEYLbzTxKtnjxj0LHpHB/1l9/yEzsRT8206tu+QSBMONRR2lPe9xnEhP9ITTeBgLuV
nSZzw3X1YIsiPZCv/oMD5W0zzexNfWswU3KgZruCYYaUaQs2/YsfYhkI9eYBBOQtmUdku8UqHDWE
zcE9RHO7mWKodDEVzoVrfIx+Hh/URa+Z4aVym+YU9QU5kQ3EtkUA47vnzRIygKlCmgRzrqnxIKJo
Y1pc/QJbAimCRpXKe/GKoRth1M/F6V8ZyQH33n0vAf/WnCIYgCaxy1+FWJj3aYZeX4KeWd+pqaI/
WNyEEZOIxQzzcQk6pGZDChN/WKE1pgPUOcLCkOuj3TaKG+3CIoTE/8Z17ODHTMYoRlbBU3PD+xVk
G/VjHK9Y9iR7qjb5s7eopGxeAA/ShffWBZ1K8fqkkT0yctoXr+JxNjmZTZE7iiSu6RaaCTW2UEc6
alSsrUlSjWxE59CacbAJNYRm5YotARPTXRGO1qyjIfyqUxs2Lpyq5inoi3FDalGcWANREFaIZNPW
7we2jWNKE5Ok/dYIGtRhjdl+/DcLzOAfvgqRS9rI6yN/5gBuuyAWo+3Nx5dNrDnsidRxJi6/H9Na
6wpyLbwjZ02XN+gONDn4zBA16S33PrwxuhIVj39wQg+F93B7E9dt+3EfUTbtL6DeeA0MB1coJuOr
7EqU1BrReMUXxZQNCcrus3ev5Dj7Apydv99qlYXF9DRog/5oIP8YqKUoDqJENejGPgiPAjBwv35R
r1mmQjvBecDpOsbcBVpsVGtPuQo0XGnV2e8CQfHxoM/54gKyHxyVRXOhtf8XzpNOhcUSm2o5IR5s
Q7kc2by+AuKXfgGkS1rNCCQP3Xpbich4D650nxK7QLcTsKI0lEpPgSrlNuF2Q9timAVnEK3fosI4
3id4x6p6dLhZ2iGrrnqxapsZ1Y3IqvuOdnil8cCm0VH9pcXCqOZz9B+h7U5nsq+5WMnQEWbFQm28
YWmQrebUkOWPjDvfzPyvp0/KweMf+1b0CL70TdkiVdU93j3raiNUgW1GYj728oZmhbtkBK9UNu4e
8p08tWi0iarphGQkIXiXSlh7lqJRBdl1qrccHytB0Y+vf1H4N10SkoOZgZqAn2ZPjUT/ciGtMhmm
HUrR5nngcMuSWB/VBa2dKs79iydtNZ2vbpCkMJJD9NA8HqmLp1lLlpXEPz1qDhE0Y5je1UjFXjpJ
Wpd14MmqvzjX+kZK2b5dk2gjTGl+ZXaWm5ZfECitYGHza41I06Ikg6cSOmifNIoPkbtGtU7pPSIX
3NwkAjLgep3W2ESAiBHgY7qZDr8GSvAOZQyejbuV0gNpmjwZadtHNZd2V1yNVPXGSbHklsesJDAY
drOf2xdhNSCXiTwstK4Kb40W8s3C92XPvFG58FmOVq28WeZhgHJBinU93bsxQhKRVnOSrQlc9zh5
5c5xbaCp2xlb7HGXGXl1J2eifxqz3IUSCavQwYmuZKphLuwHvOdqU7iApeOUvnVBGklcgmEdo7wd
Kz1tMjdHyKdxAuSNaBRBeuaLulWhDxYgw2Vf06UU1/qnLph13qoc6TVgzsADWl5X/2/Uys1ClXiW
R59Poa8aYnuzwcbOeuTLW9bMoiFJHK1mcd5vO3wJQrkRMwjcjFNDu5g7JQXavsu7iTSImQ+JMref
HYg1V9HSMW8FR13ysN4tbvI0JdtJaXUQXmSKDdLGT/QU+lPkUEawYvyLjL3WtqAveu1kI7tVVZ8d
D/qzRJg6VecatPsi+SNEXiq9R5TVn5pQSiCmMXklxspwauHIMnHeQxpy+9TUwwBSlB70Hhxly2gP
wr8qJZYj80N7KdpBM/ypOh3H36eDZi5i+cgo5l4Yiv3qFKXAvnZvb56KRmNlJkmbuMFCuuPCOI7o
OSXuDn7Tf2awCtcn5Agl9iVjpRS8/h3dmVvumWSiLUJ7VOttLAEEHxS2aR46dm2KV83ch+ACRdqT
R6h8olyPVmeeL29Ipzz4HgWU7UBujR86ffQH2N0+R68+g8mDUyDzd4fS+95q776XCxveIiR+7nfw
xvapl8oSQqtxui/HhCuFJo+bGvTFQ5mvKvQr7ELGABRJW/K0t4GiNwhAd04yR4vQX6K9W/JuQOLv
o02Gy723IOmrgirhpo5zhfV1cMolzP6ws4gokivxJBa9kuKkcDKGoYQM1ZISmwXviWMNRNZr6yan
KbJgWDBV998pQ6wtguaOuKoIi3ndGJ5Mhd3mPoj7iIww5gltLJTS7MVAt1hSCDDzs6kihHnzMsQW
/BclmFw63ZVHU4Eqg0n/T8YXwmlMWuwMxrRaXWu52IbnbEI2pZKoORCCF7M07+1lHyv9hVWSMDgp
bfocjTqDVFuvUh7EsJBe6NDWRepBuLikpTCW5oaZJfbXQQfgPXkGgd4OaXEYWyCOVSrG87BkbKdm
REzLc9WyGa+UkzmtJRa1rvn5CP9oh9BUuXbaTvc/hN68lPBoyZeFOZn2uNASiJlrruZ1t8FDvhLu
9SBWPbYHyl3Khn8BITBbKHzMcdYSURHB9wYp6z5pbgU8Cj64SbkH7W0X9EMLIfkqFY7G+YEooe/B
2Wf6I1ZDYG8sRWLjGoAwfTTm61/Jf7mSIUNVT/0vqe2bUETnQQNK3t3gVpjfKmep4rzjY5RalYu5
LHyx0d+CymVvNrUNHLTvUoscVtwtQCesswEbwH11/xtWt1crc4Tn9A4GiBasjsVxBzQsa9k/pp9o
W1TxQhzCtM8x0TIW6JTTnEMe3Clq/9L1PWpfmD7ccx9ChVwY0CmmI4RUoODSZ/xT8jIP1cbLEyKZ
1nClREiwa6wlRS+gmx7M78tEhD04I1v/PeRcW8oADt46ZxIFa9aTgfgWFFzExDqPbk6m2uz1flt/
4IVC+AIzoZLrIVU/7oCB1GZRf2cnHhvy6hn5ffcFrDDk0hVRdaZIk5V1KhIb5gV/04OtPO3KrWko
m0bLLMSFTA9IhBaXI0n17GNGRySLv1nb2yTfG3o//DPP85qRffHjL4yBDpndth1CBTspJcJ1kOx5
SW3uzCR/EzJI0D8mA0MtBEnNmFmkefwG1OpQgUrG0xN9n3DSwBAnYD2InM5H6O1DJ9SnCicaJsFW
mlYPz65XftPBhosHjR1yAUKmHPQszhEm/eZW0jUVLkhollyndHILK71CdrEZNswa0TXGESk2hIG8
YH1JYIDu8IuYsj1NHl79TV23xWIBl6fuPSjwf3lWXfQjd8AWfQ+BTSwguZQXVoNQCES5vbJCo0+N
RVLiQSFwsRaeeAzDWvyRNyjLW26bFlf4E6WSwjvUCDl4w4P6ysicyoYewDec3wyioIOoEXcYnJ/9
wNSsv+61FmnWmWnD3DrUVwElWZo57JvM0FlTw7FMuIEyY96AF09U2aL9TTxafhFujV0M1cyeiJLn
eZukVsmuDAMzO9COiFj2kfHvgV+Nu1qRxAYxIxNl1ktReLTKZ/CaDm8aqlk1vtrNHiQqSHpE2kJL
8y12JPs8V40dggGbKzqY993/uSKigsGU9pDfP0tp4RV9Bvsc0a94ekHep53gsM8qqJLqJQOtGobG
CS8gQEVnrljJkLjuXR7MIGeX2LSchkYQpNo8j562+x/a6MMDBeBC6fNpyglNWMbSFZDDlgIoV6aA
S9NdEZ/exVfRkKTeg0taKEdqan+bDAmYsaRtmvII5eXs4XnCiu6OI3btZ8cf/CzNSXXAeOfJ8B9E
68iEwlXbUcXlWJhQAqCmbPgQtqfpaCD4yxmiqoBmaxV3JiKdTh6p5o6Qr6u+OPwF6YFDEITCTZaK
RSvNCpTfRfEYCVFGpgvwYL2NS13VnLWO35H1t83G7vSVt6MXu/otFHbjvTQ+yfGUzkGH2PZDK05J
idI9tL/RRRR91aSDUjPZv4ICnQxqrpHZqTdF2AeD6m6XPOY0cnRiocOk0LlpHeJwtKRnNkoARFnb
gqNxxPNXERTntSoPm4gDYvRalLGKfq8wEcHKX62mA9poR/bT2/EpDMwMpJoC5rjKBN1CyvEw9gFK
SegrE6tc20KDgYKbQBaX6RfHOzr9Z1Hs5bNVikLwY6J7iawlXZLYElw0YHWZD7nBxZjy5ufS6lCa
I6bMIYA76gsjtYXwKQV4YmJrnlyqoVitj+xsXzqIT7jCeqGHzWOcyLW6WSXmMEw50WrCXiqVkjxc
2RYG8hqlTDblEL/hFaHf84gpZWR5piK9cszHBvWQsk95JHR1yKg5J1enHmJLSquU9ON2ArMeg8/z
6RNCrcWdvRvYIzduUBCMEnSd9EmTWNEjZqmJ2zUwFzrS57QaGXVLDX/g9GH+TRcWC3Im7op38i5f
HY7rUfRT8jG7zmyz7ZlPOReEvaFBQStHiRnLw17aTAqlAMHwQBy0gJaCjRIMqR3SfYupsvEWt8Fz
VnJb4Pc++da2+aD7lfyjs/3YYRihbUlbalkxjAwvwTAqlhjXmeZvOCz0PH06g+QJMYyF/OmpYbmR
cq4w9RlpgfLJaUUXFujD6bUsfBKQJPoMAROqQYDd6WzpIt5OA4nuBeVJHO1y+J7xVAaglNs6zrbG
TXxMoZ956mnLg4N9etJ0UI/2xf0i4j2AbEmh7wfwODXg/bdNJS9pkLLMMmWL7Zl3ygb0gOY9yvAy
jq/olXTZ2Oy8bmGEkuln4E1uOMlll0SZQJS7AOYJZy1E25uK/DxAwmivn/k1FqSxQB1k/1sck9y/
64EukRGQbqR3eeAxRLrP/nwjAO0r756vcoCUXxFTkeqCWrNwHrnkOglhQdG9M9uQEqQ04VWOed6d
dhCiWTrm/WBFjHLASyFdqQq+zUpSrDagcgfemAWonE1KGXKQ7T/70QI+KPU1YlpftTG+HVhqh/qH
mCCJcfoYmEjTGM7yej1bq2UOe7iWdOermlKndzUVzsv2QDkNdQsRA/jK+JQknklQ8sNhiVhea4VZ
ZgdTHX/5OZjSMrg+rwwwuXZ2tDnGPqoSfovV1Kr8x2JerQw3rl3CxNWlakmOZmYyNnboJxCzFTBO
LTljIcL+COinnfvlb2arnMWoR5nUScyMuEbrxjexR8I7+GyhsrdqCyz1/9ZPlRIQ+jFZYq2aOHSt
oyCGcfXpGL6Q1CGbAKeeUSh8hcXoIdhv9cAurgRMkvDr86F9kuZjn3eaulX624zCj4UVfLIAuuSQ
LdGIoIagQdTDYdrdFm0mpldGr1UNWAp+pXWrxc65svDbim3o8L4CRN/TyI79DVlaZlocAs7JAihu
SGYv8E+QRwxgHLHVN/cwJULI5AqeoZv9dZuY9dZyMXdJ9ss+kfaDAdOJnTNHvt9LCQzoBcB5M569
1K7F2dhy7wxeaBpGNmb+87dznY/M2GcpumK7vnRNdmDdYMwUGW4T/0V4KE6QOOFJy8aZRGax6qxC
eHuZcY2ImW4pY4l4Q3m8StuTqEDFabAtuMQge1ORJOAZmItUZcJRYqLHylghU7DbSmMqWZNK5UFU
I7oq9Dd4P6l5F7yaZP3gygebWmQUJwEOcdJhWMayFP2MSFMCp6TR03IfRB8MiEKpK3POvXo0MPII
dLKt0PmlguldPlatDJHqSjMheViCd42nueCO2Bj4QfdTnjuB7yop5FSjwAX/JYS+Q01b+Y6r5mcw
XoTsSs1htU1pXInM0cKlpdrEXBitvDQ7InmH8sAsvjJgfE8+Lke9w9tE6BYpYtVuExulEL0s/fLj
eiMK5NZz3/MSJu4RteVksVqvfZtW8rT3d/5826LqYdMHuV9Npp31xfBNlvq36OmKaTEFhluiKVRW
/7Tv1KhEuIWMDO7t4AA4Hvp1V189jE1IQTtMq8/2BUdZlPFZIqaryYdwMDp6ilTrUhiLypniSNvZ
xWKyADBnaJCoWyDOB8ruYy7hG65aWbD/CqroGAts13kqzemQ8tNKa/dwOuUG1/Hws8sp0Ut9yLvK
vywgjyqwqm4UWWd5F5c1HOS8dQF2HI4Xxs0FxkQUf/uxwwN/oBoxcENeiBxZ0wzTIpehj0IUHmd9
z9oRt5HZTKCVxOX84NctBS66YazZzEAcBxZRRM6YCYfxH2MxD3sbZwzOhf3FYBs82SVZTXjD0MUn
v5OZpU9o5RAgrGHrVtFdcTVMnMj/E4pRzORQIGVP6m1hOBHkBubk4JuxSmIh2FxlgEMEynzoT4z8
6wtbu3lnwEcg6mQ29dVor4h96BQUT7zPOmGmg13UJqQ2bwVJI25qb4JVuOB0iXMEJBW41P5YAQc9
PqQ0LLF0QaOarMIthf6eiA5T1XgbSySXsCnzgTL24eaofLQsR+BZwXpZvwGtET89heXEqR0n0qqj
TfAzrAnOePytUe3+vNfsutep7IMDAGXIRYoo54kssL+B4XOhbhXpiBnppIPhYNdUSGWYnl1ZtO4w
WGPzDl5RLbAnITrXw91r5MEEClENa1C4eR70dUVURx0Nr/C2Db+nJ4a6o6Ej0i/cqZqR7Gi94OEl
uoogUrdEOmZauq4qAanCYehdjMLtM8YnkQHeCHL2aA4g7EXUWM91pILqr/ief7gCUSvFX+O3I4FN
m+mG8x57z6PqJHl6BGJN8VbhBvf4h+J0xL/ty8vELdok5ZWQEXXl/vLc0ijW39XXlzeePhVY9BYC
czyLtG8NkontHriUUwLh5B+xHVYYA7txOUeZds8ubgow3Xiwv+GbKI05WetbZea1dPXRkx482CjB
SoarP0FzQ637V2nQfeX34th4FDQgUgXhBwSh2S9gUo6sfWpZSATIEqu9xYxZdGgvkxeZ1zBbalFn
XvqVTsxu1K8gzau33XqHgoxTOTTGkqAfBZ5JyZX/Tahe+EVE8I5iJUTiomA2jR3Y/XtvtrloKtpQ
Bvid4Mph7RIsDh7QdWgROcYXEDcJyQ5qj8Pf80xwgd26scD13FJ9tmQdgSlQnfKplvAnupBw4VEr
25CIoDkRbtBKDOEJUtrBkuCqLFmfV127lb/O4AGLwPdeLPhU0KBnRCCl9WGd1O1kdC+czDxFJI9z
WDNxtewbROfZ1miDtcEeQp9Lbk4LnUI5B/bd5AKDgydt5lAXgxrsSzXid4YXiVmQSRHPmTgt2tQP
1E47kV5nv8e4LL4V55upLIMqJdcNS73COlbJCX4CqlUHmddmXH+jW+AW83ccX+WD2loUcT0smXPa
gf4vH3h+jiwrPeoRTrV2sVrkUpd/AKlx8ttjwoUEFWjKJFMJfYd/Z/h/AheIMOyzsKeNy/hUUcwd
NPd+l6mswMcWFtvrPlqte/lWXtmeS224IbChbqNgFJRMfrBsw10o/02+6rFOPmCIauyKVdvl5I94
/IRIgquXjfozEFpT/k5sGIs/GzUK1SuGXwzjyfWk0juvaYAdqCTaETL0JGPoDp7fsGt+XFrawKcm
4Rory0YU1FY0QDeA56QA/r/9YeD1I2HHUOYKZmjuJg7T73rpjXMAnjQ+e75mTlpSjMT0HUs+J+uM
3YqR2Gfyz9VB5LjJrxYRxLOb0z59QuE4kTMiHu4ItJH5L++9Br34Kd7V0mA9G1RO7ytvsjkxR6Ot
630aS5TVSH/S0lEL3sM6GoUQpL0+XeR0VVgvJgBOntqLI/9IVZedX4Sn0TzfjEV3HW1EKaS0E1X6
qS4DGpOUaqJqqAkuVhXnLYHKLsgkOV+HBNE8fta+ngDp6KU/3QdmcLkOm2dPsy1PIgtGpTeUbLl5
vMBr0V+J4gjLkVtqyagSZiOGiEmN/Smz83esNSb2VcCBS6f0I/hkGe+mX5ebyGi1D+rPdrBazhxS
jORq28Eij5rtqEEPYBZQF5vicD+joCc5+i3P2kZd0ncfzPOdYBrWsP7022lZACSxSPqXWJqNXGkk
uGAJRBa3h7jTvp3aeNWJVe9SRBRCqllXGdGm833CZrm3N/VLZbwSZn7hECDkAW9SoSYxk0GH7gGJ
dRLfuJIE0RPu1nwRBzE16WYzgBbayFMKnhL3zcrbBRBd5Jxp4DHDHiNIbp9TmLZoEM5IGhC6d1g3
ozoEtwX+4vEmAMKtUsv1cYQmuJQsk80MCLnn9xJN/qDP0IdwkYJaSdo1udymXievQfDlKihZhz1h
VbumvxCIMt3jGw8UFzANr0W+NfzBuxmeSDi++kOPcqOhFOM7za4LpCmJfBzJ+4zt1YPRWG1qMa10
oXOl8oIhcoxvI58/dLS/N6JTy5wsaRXnkiI7Eqd6EVtFOgbzp77M4JrXvgNNHsCYOcjJBqBORQZZ
jcRdgw6xN8ppMoujQA8xIH7Uj71vMGynp51sCsUDVgYEFgWRUZEKShcyNaJSov+rCNsCmprXx9WD
TR5QTCvy2o9OA/nCLG4+VqfHiQBgyGdb+DtHRtZ9RpGOvp+hAAlk3yPHM2Q9LoiAVtlDnrZcRi2v
iiapY0CGeitLhQ9wjGxTZwMIxfrGx04d3aPjc9TonRDWer+khp6cosKCDLtR4hqrI1aSnBEZEba5
KPgoudukNbivVPGhvQ2PZeQZ+qhpITHNOMZ+p2/LtJirjMhuy+2KZHZ4qyFsdAGDs3HRTmGrNQ82
shxKjAkac0aAKTQREAEeOxz6TvE2ATtDkMiwzJTBAmpaHuUVcyUo4lGXfjxYkpiyqK6Ytu8kEe9S
iuL3Vs/W+vaZfVOCmCK9wu5AhmgTTyTuXud/u9pQZR1IpMem8bQA3T42HdBUKZh8kvuExCYADPBb
q9jXugixHPyOw9UiDFd8/y7PFL9//vn20V8k2G/vAgguA64girbFNfoiN2b1u69VpQSeIQz6LrTF
Y9pPLHv/dhtbH/7Aq0ix1WBKApopbxb2dAYi5Ux8gKKPP6ToPvU12FHsE/waSOjRb67N6WcoyYr7
hv3NLqoEiKXw3Fsq/tFNJhZyQzUSG7tsYSgVe/Tak+oO8cVy8ZfLfP5Rw/LsMJE2OFfSA1bSXw36
BQyFl49596EXOW75lMmsxSyMYffKjlcj8iNiIVWG9vMZtQJ+HFydWNdhQ+7u8NXpS+HssLGHoFzK
2Mwmtcu2ENxIudJPETxw4bAwx2S8algnJo7B8KfiLBkPwf73vH2iX5hmliywM2v5Flgd2CSpNtsl
iLI7g7OvuM/a+rwb1/t7w8MPKGcIFNo1T2PTHZH9R3XCrMoXVeppcl5NscYACjvgoREvIsUtIlFM
7PmkTWQ8FKab+lBYoHE6BZ4Bp1GEYAB1f5hNUwq+4RpcLScGM0NRDc6aIvia/+F6OfCfAx33MzsS
JJw2nHrZW2uNOXyH39GOi7QD8P/E9Yyaf42JyrKy+aLeQkhmnRQft+yi1j+GklXSAvl25YrUiJbH
qWlmLB3ct/xxnteJT1t57P/472rmMK9HBSKKUMxlrLorYqaUQWEzBpJxX4JeIkGoDWuvEX2k9SK6
X/4QOufo03Kq/vLDX7Cr6gP2sN+kH5mNOMC8AlgSw53ulRJDjpV4DMF2ISzRIS3SPTuMMbdDU8nW
zHnIoojnLp12wd5/bz1Nrktoyco2Hi5exnrTsTd0H5Ih0C6lNPqYzjZ/2lMTxYTwtTdwRRlIwI0t
V351G0OIvuFKMjCJIlRS2rycmfMlA7+0xIhAEaEJq5HfPi/C99dBaSFWyx78lezD3pwCHZCm6New
LvHlFqgujDW8qJmfX1Hx2PRThbfre4Pbo2iqTO5J05IOKh/eZRZVihtIJoNfm3HOy9R8dr2iV3DS
Zhhe07E7/574QUQxXNa6nIAh7W24EsgOnfuUxy4mA75CfJD5rVBwANz1F1m76fiupQypVRiqGlQo
pdVLBKy0iGCxoIzI46hkVC+k7uE9VYJ1l+NplUor0hM+WepM02ES7CkPZ1s3ENfBDmiU3PxEVttl
xOEHN1/8o1QwLDlKpJ2opug9sh2MLV6FmruJ28lA6BTg/6QcqCW+7CTwaXu84aDWX7kV4xDWWcZ9
KsXJVuZYzXkp3+4yjn+BzE/HrsntVj+5TsGdCghQxozeOL6/YG7+k5H9FX5Cz0sry34sc67sdFXp
h47i7xuHwI+KDR/G1bf3Aa7XDmjXMjmG6eq/2kYNvvWe77xnnM7WAJCGtYxw/K3JjVe1SOoaYj2l
GBybX6avGgexfXDsd3dXOBeJNyfIyV/a2DV00vhqAvdIzKQHjq8Lp+sp0gpE/+Zxpt25DwHM0LmS
sbgYY8H4T7g0xG/wl1TUCUYXO3d/utv7I4A+K5l9rW8KdPyY+Q7tULi/9F6to8XMHYyQTTcPT49O
LBlkaafIwPKpeTVwoSfXoPBoTrIwlA/t9WMC+HiWEZLP6hJ/30A+sOmhyvs6tPu6ci43V0bC4sWj
W+U711ivU2pBVSz8g2AFh/xDvvdeC3ZgnbOfqmtlz4auzlx9MVsc08IkKVJZ22nZoY/qODTvbl4k
XYH+bc531eK7Ht6c415cJy1H8I5lSrNmbH8UwtGhm7OYm30jUHPKCNc2Hx347mgcFoa4WZ9IhxAT
sdYTvAGG8GTomzGgEcZRE72cvSJ307bIQVaOKne5H7vZAsuSElS+A4Ihk4AIZjLvsxePYoX0+wpb
rZw3DUoJzZ+7s4ZvkaSm2pOgb9a7lYV5zNymYEFRWtNiqt+Ef+4TZxAdK0/mbLr4t1eMdKK0O/Cu
KMTpumuObbwzE8WHh6q/2WbsJEkwWrBfmwYdC8erTwiExQhBgd+Fd8ES56cpb5dkO7wPowLP+v08
njmZY1V/Y0ZIuEmJT+lxmUxxtlEkzJcJGuBZLQkYHPrs1Foxs+VF4woBW2yKWM0TsTsRmdUB+6C5
zreWmseCD85PhIhOolOxIDQbxNs2yMysTgaoDP8BZaRYPOyZJmNIlffctLs3N8kQlk2o5Pyl92y4
5MhphVMJhrAxh6W6TnUZG9rEA7Y0Bmpx+jakOLaIZvNTRaLYh1i9ubRj00GkGZ5amEjN0FEatbyy
iytpV+TWGe+WQZL3T7IDvzOsJ32GcuVtAiVUsQ3Dk1emFMzJcwcF9g9AIgm/u9ndiU4rIVFotV9v
VBtAIAMzu3Ada+Rwm6Fl81e90fU6DLb4y5l4diAapJOFAVnvpoUou1c+dXpe3Kko1BVeTp3qeTD3
/n48nn/YolKWJaj4JnbH8NpWnOTJaR31spQhVxP7ERixloovtldSbfE9dyUZRfxh5DAXJljKB62k
rBzqvYWrbyRAuv2UWFdMbjfb9OWn5w8V9SPtAtvu/gCTfeEm/hVJ3vcm90KaV0wbvR8xz4ST6MhZ
dKutPN5m15Sul+st/kuU2vSLLBwMhBhDMWWxLB9fygI4aakz8cRIs12QFYnXCW9e0O8MNM9NV9Vq
V2QQJQNOP5cw6fcGKgZKdu05P9ahWVK79zL5uCxaW0Ld1jGR4KklT6xBLRpKRgeNi59I82vLr9cM
yZgVLPu3dm01JBzaXJdPXSzFg9UkImG/v7dvWQUh4Ql3ddDazCVYiVTmEumrMdJFu+jLFpcTO2OI
fqfsJsLH0RiEr1Gnxjtz+aab9P1hL6yAY95gQ1G2P09wO5pG5T563ISM/am8vNyXUlaWUrELc3+Q
e/C6B+NYsR3fzDtHC+8LITxHD2FK7Mkkw5r+yy6/LUoR4m83YNEvXBwWE+e8rkYoFa+wjSxdhE9T
4KiMzmiL76i4E99cQzxdew6gUoTllU+5M8vi5NPIClBvBIqQBEmvD+NTM/LySmV9CQYp5yv7HK1A
I7F52UfoC8VRCRKBH95arfAZEsSm8akFBjoWRYrc6xe3La72PbWL0/kKMrEMi6qFfIyh4PuI2UDo
zCYyTUomCfKTtaMFMk6B1eJkUoA0IaIGXdxoFsCjhTo4tzt0Xztu3yx3NfBNtQ2uiCp6agnCsjQu
ve2f25IUrbAbm2AEZiczSYfhxXPaZSRHHdzMx8FU7HvvKoxmnMqplnkswVKJqr5lC9lw38tW7loR
DsftOxGRg23FNgYuAWvM5h0Z5wxMW0/u3+LGJj75c4bn+bQfBP0PC1BhwQEt4RBtzhD8xpwJQYiE
5Z7ldh71feEAUQfOrqhu7NBdPZY9lUU98TYPvqa1dPKYI8fLkBfo0rNMhcU6uyhNBWLRNhhoD8UW
PIGiPuChDj8j+6vs0k3vZiFYYKassqM6kV7KiWpp+ihNpUMCSh1zIwq3HxP/U54DuXfjKiaaX3ab
7kF5NHCkIOH0VEX9ykuMF+0lYlSajgfA/gdZClRGArimX1AsnyGOg9wZchnOsh8Hx4sQW6Whi1dc
YwnmSouz5i8GnnX1NeqJXBIXzvB6rouSt1N8/ekDGjtFhYwhv+466sXDKGGSc7kzvm+twD7P5p48
53NZIvpGTgOOdKZ0dsT6JxC2LGwPLzPCQcRiXipEscbM9AWaa8iUYw1By7VliNKzGKJZDD3bJvTE
B1KAJBGGqgnzu5RXWi5XTCNunZyPOZDRaGNtgUymT2gahTgHJP0cYAdQYv7TCkK1SIdpxV1Zml2b
EC7Fres/SiQ41bSFqCEtLnhyWwYw/yzBfxZJuAvGY/cMVGcmvETKhS+oFrevY1cc+qv5I7khd5QW
QILHfiJHWtXZSixBbXvalQiiU3oWEzmt9BL5s7KhtMvCEt3N5q36E92YH0mdgdcX1ZD6t1K9tnC7
1IvT8o7tmaw1yIpfVb4Zw296hKzn3i/ggG+lR1qgkNe/tuM9dUzrPqjvKAo3sbkSL3nGNmqs84nK
Mhne1US4YvuHAmMb1bAFkjkwf7hUcM4l6jHT9v+ZZJs3cifDGikJBtNbmda1rfC7vnpadF1xbkXn
52RIMcS3P6/8PYHQ0qLDvIAElzMmXkvF/WEOrAUEISerkjCjRy2aLjYikdIJ5a0WBFmhFdZ4llKJ
6PZ7Tc9VZ9ruLkNUv8v68wbvdwlmefLMe8WsKTJXTztDxuvKLGllDhl6vayD7aIORKyyotiAk3ry
UJc50iEOlIDw8sUl/zhzL911z2hFzRu9rEavyt4tnza5gQXPo0KAKoGTJfC8xtDgdN1ZBZAKLhhx
laOk9hinL9sz3MSyVi866VVp0FqBbrEpC/bYm4AN403ZrhhmS+mV4yHeK1XRblgDnwK1MX034ecy
2azz+H1ToUMCuE2nSR+cCO/o9gatkGukKR+QN48aMQFnE8FZvrW49HTbgEwqoLKT7uwx4qFUC/8X
iyDRcAi+fLOzXEpOrubUx1LtFDLpWzBTDpfmUJ4swvKXMM4fuVPVQN1lttbFYNN6g+ZZrY3CYQdu
5IMfR8biXt/yzxxeux3v9sOGbvc/3kbJ7A+0RYwczFkVc1U0zlxsc49qudk6mx79UX2SDLe/v8bY
wlymfmQAoaIUpcyiEnVYZ4wn8+vg3etfLfiIXOSk1WcS1yVAoXwosPgL3QeJ4o1BuPFXx5NElF3Q
t0SquYhket8R58jHVtUcRmRuQY4/asZs0skqFh7j4WFO94phMVJ1S8GngaCDd5PYclCaOdmjLfLY
cEitJIHt5FlVI1Mv1oNHll5yJ5q5kcievL/xMOeLXqTN7nSbHOXvLTtHYMwHU5ZpVAXarECIp4Qx
soilv6HZz/rZ5xoCoyH8mJMgr/4Sv0ZvjguEmVRrCFI9jlA69Ivl3qThPh0CfmCz96sPGY/jjsoX
f/AXt0AwbnU91CVDSceud7K0mbO7ZnvcUpTqFoyzJtZfNPlztaBFruDmh7jMyZdF4bromttLpQR6
rU3NqZRMJv4xCDXdsr/Ck5W/+3UmcPlkHkynlJE2+m8bCgQdL8ip32wYNBF0zCTZPx/tHgko2RYA
DbRlwCR/qQ95AAk2D242Up4SoCAIxdGwiSCzl4OumhIV1FQC6VMLyl72zQQUQIRZfnX2WDOSdt6m
mWhhu+mkfmwuR0xRNVhEKmodcDTYhfEhZ4VtdW7S3JpFX6VHeiainsVLpdDhtDnlKeA65fWJLrZS
36Z/wSYZiUNpe4kAfFoj2fR2J0nHeJRvdYmRQgW0Slzp5Ieie2J/Reqi4+yvmNbgmwCTs/Fv/Dac
Fv1IWQ5C/WiRskEz+6HblwUWZ+vLtkcABcGsSbmrDPM8J8pmiN8/HFVmSk+NgNJ2Myl1LynsHDAO
dlAiY7cqv9vG+q0DOrtIxxKI6c8py52SMmVYGRIzd95hZ1Hmk5PeuXrjJ5kaD0x76dZ1VKoYFSaR
GbnLcIGjZCoVI4GFFAl6hrIbo0020YPDIuEePWGQncpPPDigFcj0YU1NI5ePcMfBYs1/abqe0enr
VqXkdhUKAV3ZC/5Af/Y3DYWun+vCxPC0S1jJKluhSP2afv5JzZ9WMmDP9bcBLo+pGRjmxbajdUZs
kygdIJTSU4xf8U2iOavEN78qWz7xOUr8E1pOYV5aJGMniCkGRV0TttnTprMgMiDVp/GW63ErUV9H
kaKO8FNtXdrIFwNODYFt8QAojSv3nCn1JrlrbgP+gPyDTM3c/LdujbPR1BLeIXiwdM/TRxXsuzNn
YUlw8xA/7tP7fFxBAcvDv4XqSeHOP3DB3hkh1e3y3qhyBcWMRV4QwSAH67uo6Cn6PRYoiN6jukIS
Gi5+0RofRZzHboa2LV8V1lDp42dgzYHu4okUqCEtaPGSjW6F6yTxaYFHsgnKKrTDIljb+VWPEq8x
XZqvyg6JNdnIxb6n0WzVCxsL7XWXer4rlpVjWXwJGSgvVbwi8hKVlpESEGKwMbG3abxHoo+TO9IO
QWoqXad0C2n0DrxLLDOR9P6BiFeNAUupuOebTVLx1xgTrSnqffetNybVNje2Yoz6+1Bd6vN1kIAw
kvJ5mq9oC5RfkZro2f2NGrpyBFz9HVRkJv4ODnyEYvFKaUulncpZ61ubDizDaynqpB3rOCP4a7Uv
u+RevHYPWWvhQHAP1bLtsvaAK4vOzXNMGkDU80RPcfGY75bYoXur4KPh9d2oiuA2vWK2xcTLUpvq
vBRSj8MYotDR6p/UNbd4J7YWZp6GYV/Zl5r9WM3iERNAL0+JYqVo6uFgEGS7U4m7T+mQnHWqTVd2
1wetjTYFjOwqKC1jFONOS8c9jc8xLYELX+fNV1PmNfeU4fWnz5WhfxHzaV24lVacaqKNH1q1KRmC
3uzlStBK5VbAlMluASFRbUkb0EWkW3mhVWtS6WJNSq02D8U/Sj90XSRt5bthHrSS2twl7+LDCx6C
ptobbEnRH5pHvQ6Mrjgbs4oo5yeWv8s4R6afLi7Fa9vkNhLeM2PDg2nO+r4/RwGMXpFzglx5QR9v
OQoZrWUxmVf0MnaZbiKvQq6Cb6MXq/xcHd85oHwYW3Iymr0fil+SK8sQqCi7qjBX9hYKm7mnWSnx
Q6sIcJ4z7f7dYKmzM/4jZI6p+xdfeT8ZvWtLNmI1ekQ+Sa8C69s30VfdUIeXaCR60i3R7V/vUeiZ
kpZoMfkElweE/wSu1dcn/Nl27NNG6xvGl+GtxI73NPJZ3O3qFCHJj50zHQ4UuiRIW6bgJUSDtzuS
6xNqFhBDGnxqZ1+fPensW5b+OYAu+l9teb4GiK+22FqjtWuLxX5AeuQjxS3UIE8ItE7cnWcAC74n
MqudF4Ab3ZhuulPqITjCZy7GtB00k/QaIQpRCQfQqiMaK1t1G25qx43iQHSOdR8Ygc2BDFicmTAE
/fPEzNhQFM6s8tnmg3qTKyTl//N1ArhXH04JTYPfkwk+5S6bmVqTEFJaBaL3GLzrFTlmKOhkuzPr
kCIu7Bvfl+7h9NDtJe3KAqZaYCtCxaZH7lfjnfPExHuuHN2iwiMgT+5/JXJ9rayQ3rKfDy6KQlQz
W09/aPh542OTiV56mGxDV7GtHYGI7pmWSKLQrd7el3Yg/NO0IQPsR/l7tifB6uA5LrQ4MsURZC5J
kugZ1qkpKgki26k39xxPZJagv33Tnq/FmrrzWhztKf3qh0SfhEeibHiHL8JjVBlWwWd3kw+KbK1D
xcjjWaSaRm2QYolDRL5XguLi/CYj+yWuWJH0EWWkCI26ciG/je3171MI0KeB2N3yuMOHF3lvY0lK
4+7jOx1mNPJQSvZL27IvnYJ6ldSJx5pSMGImFtYh+HaWKH1Rw68VuqHUALeRtBtdYMatoVFpPlxj
wXHi9BqpCKzfJM4jckPYbl/gSy4AtdYdGQZPnKQZlT+34GAFV9drbR3aHulEKPSsgRDrdi286WjT
DYBDf129p27E7DGI2RGejDTN4nDOZhBEBVEENwUCUAs66f8bzt24B8WejlHjhf/w0SPt6VKlTacX
Vj4Jb7RHdp/95AL/PHFPdzIkrJHh/UvtnIYFB96K80k6csPIXlvMge1SrW03qDtungxLC8fCC9jM
ZwafLNM5HeED3eVTeoeOkBbwWuhuTuxmI+5NjMkU+AL7uTCIuhGpOPuBFH79Rosm/yI4u5OKOCTv
2WcwA0kM9CU2cc3NT+HfauwiU8Qm1y413rhzq96tg2s1pYGbWkJZmeTydDJqdeaVIhITclh1aD7+
mK5xxfMo1H94LeIaMuThHkxYYfCwI20Vr+/S6+N7bKfYRLWKoXx5weqS6CLTIokF2nEztuDyfMer
J69zG2Pg9NNV6yWxO3yVoMDEbGUJFYCguoXSH0UW2mPirV6C8qHWv4mBrtmNkFJW4ULnXEIGl+bZ
XBLWM/rg8dEIBMUn/vRB8mG4fmgzlK58Bhy1McgBIu5sCj1D2Xk/KF0AJ3duN0IvGhZOnxMC5e2X
0BvSy/odqXPnF8HFIgwW5MJG6fu2gEzybimKqRKrYL1qRZIckethXkOFshlYn3Po9g1A8XrkpSvS
6esjJlH4cwdcOqrncPG1C4xuDxg8DtFPFNg6/y1miQvcqLO2Acr3XEsafGeVJNPSNs3S4MjBj0lh
NM8SP14YuEJrtS/vjY7FLn52xai+RsMDjEk5WQXpJcbP4KG4ocGiwKs7g5qbryJ9s6/dkOz30B8m
t3rHK3MMsIC8n+q1RDz5mBP/5q1NEUnOHkxSikI9yu28nx3JciNQ71XN/JRVITlHGHJDw2LdPLHA
YSFLF7G8De6rmaUIufFDTG2AUBrKY3YLtlarXsvalQm9CzdCrbLeIk0nNWIF2aBsVbKFNEM/ntW0
ONO/De+MkdJsGSU+/8YOldTrhreLmKDK/GBPMRdD3oTQ36ocEVzoc70AtNqee5LtFAmmn+M2+/V7
Y75Z0+miCBoy09udQikPWp1rVSdnSUzEJx4pB4a72lOd0lzNYgkXtjAiMumHOvBgK05u4FiVpwpf
MBOV4F3vXI01k4cB9libFrR+K8K5J3BhZgM8cqPAm1556rYaQpGcSftxHGWN4FpwH0hCNzVkGtAi
QM/CZX4ERut8c++81P1DDS//EUAUnn1+LgE/+2I/94P09gI5Q4WD0DvKUVdflAHfMpisDbhC/DT3
8ZmNCDU9w7jqYwSiI+fK1HMWJWSRfSmEMXK3CWTCjDfog1k4oxXNKJS/NKVeZFjOMOtkJErEI6JZ
G3l0pDXQFlgWnDiQFgtmNXxL5hQSOOSir4UhyaTc8eH0zC1c3LeRsumq4knnciix8LKET619VCAU
iHdCPXjcltx6UmwAKLhhjoEIGrug/AXlU68G1xm2LjzxcMYDyxm1EFX/L2AgmEY9UxfGBZdHXPvz
2I5PT1A+/TkOGl66Iner6USomw6HTfg5F2+PoPTEf0Z2NoUcDhNEGkmxTiMcm90RGg43jiYrHVzB
iVO+jziUDbmn6vdevco9PJsdkOzKWLif7xFuo5TRC4HdGWCwstIuImJtkg6jPn+5O1nLIl+0B8Dk
gLxdZL5Lx6u0ORtKTnfjN+W1gV4b6slc3Qe6NaXIjIr21SGs6gQCXJMc3VqUikzD5DKQgCu4FMiF
7YAAXLQ9daV4Gs6YN1PqaJn9t6sJ9dozbFJmMIC/sH2nLiCnjvg+qQaUntY0zEhPmVgPz8nzjkl2
vuRdQ5l0fFkBybAETDMbrLKhpRPWJ3kN9Bi+qTKUpM9Vn4ym9qhIs0sI+UJir4a86Vt5ZfOTPDH/
OYQEWj/vi7tmrYcXc2cSCLtlnffXb/GCYXn6cATzgEa+wdzz/bm2B6oKkcyy0Ip+wQtBIh/s+aTI
oMmV3KO5atVQGTVSkNEfslMy1j0wzJuIya0brg6z/R34bnIEVk9222dD7I52vdTMQytpynm24RO/
2nfLybsbf5RgNs0SxOh8I1NxHTckAG29vppREKHv15CTa2xlwg9T/ocXviRIER4naumFBkU+12vC
nnUvUWCpbkLJ8Z84Ze9m7deVEGdMjTDB0MG7lME4RzTtSFMRqgrq2lL6Dz+zQz6pTZJ2RSkahi9h
qAMPrCqc+nrLT8OpidDQSklMegDfppK9vc5NsYcmETlk/hZDRMv9yUA4Fmfsh71hmRZNVuF54uXf
VZuWFX8qJkS57AxkSXlczZQGN0EG8yJ0WhkaA5dmoYXH5i/apFLEmM0PqTy/Oh1HdsvNkq64d5Gb
ulZv0tOkFZrpRpaJp9YpCuEwiLPTGOwSTPVPr2ZPos8Cuhnpy2W26cfSeBlv/cRz81A7tRQF0XFa
tWSThhmhWAOT0v8lPStlBmQ3ZaR1fUgd+hegnNq0U40eQnQt4s18vcYCmWddWeJg0uC4FsCLoCVs
fbmseA6uz/HXAs6jLHzBsGj8NgCCdLIsu6xqjGev7TUYre/ozwW4Lu2hf6TDtZ64MtcfHQ8HbBf0
3zCX29kBqaqkBrUuFZv8OpUSSH3TTMvtEheXo/OeV4NOxndte0Bwvu5nH8/mBVvV8SZqJhK2E0CU
x6YNSm0eDkNq6H/mjTgtU2WSTQ48dFw1cMVmZ70kmitYeaBnHKJO+HodIw7v3R0DPjCRwYIG8jjH
iGJ+zZOeGrmUD0ErPOig4yemoRhrkeAuOtN/w0bzR/3NKGrXCE1QfjMK0S/xUDh5XGhpSXKUD2BD
AygFophaficq27ZLUcDldBX98T+pASV+KpdAeCu5wjOwMT+lUYYRxUk7linEfOycJB0SqsqlemfC
y8AJmxP7DYRYeoIu4RnGK8sYM/ygJg06i8/lW/SlZAv6jNfTxUfzE1hqt2ZdCUt7BOk0NF1aloks
2HBEjMRvpyFEqjQci1DdW1ycefxuAIk6Irl0Ee3VezVeP9wbVDZmKzjZ51Fm47YlYcvWSGmmKTgT
qIATceIvbYJo5pOuLceI7Km/i3hgzax4UclRNDMsZnRIZdw3Asu1M50iE9tRVSr56XGkeZAbBD6S
yz784xki/S026g/gqFVnvNePP+X1NygBd5hHrDnUyU/boGkeHJPnBv/kvWXLu4hSagItwMhxBmXs
YnfYWqEEVViCxKZkVtit5QQWpi7L/dPLjkALvKHRCJYMVjtnFJefqG143cub0UCQMByc6Yc2vhOC
4BibleLS/+yC12U7FwjHsCquuEPHKIsWUo/CeKOg+u1iW9gRJWH4g35ujDPHn3WWY6o4V/PSpZwA
02FVkxhTkGugA9eM5LQAEtTkmogL8EaH2kG7JHZK1SSI0u1MLu1LzpWG+XvHNvk/kvcAKNuGf/V5
zXtmmL5pnNvKN/QshbLE83vtVzxuani2fP00CigWN6EB8/rP50KKYLYxgeUAu05A4zcSOrYRlmdL
hG3T9dYd0Pny7EiCfXypVEg8mw9n9o9hI67mkv7kglItXGaO0DnDG1Iuc+h4QlIU/Fnm5WoXPZBW
SRXN/apPZJfCEZMS5rguffc8pLbu8XMbA6svHmL3CssTAq1A+Xf+l/dQfLo9hztaPXas3DaqK8X+
HlXX18j9TV9yrXRBlXQrZLdCm9p8fFu3L5ysEcuh5bEQKi7uIISu54pXwL/FXGS6qwYrPmfL1DZ6
n2CJ0wuj41tENATeTBVuE7v0Nxr/9on2KfL1GCcHeru8zK8/n19nUpg7KPbFkK+BfsGoJiAW2QA+
e2SLgPVox3CEVvwvVf8Zpb55WQf4/ch1kTXvuEzP6sMEM2toQT10xVrZcmL9yhFDdltM2rwz+O0G
1zOf/bumXFZHWe4rQ/exQCXvziaoyGs4DqNR2/+LZknMpuZ+4CH17FsJAslJ8LkY/c7QzFwCbno4
P1BHCn+PXSr5cIufrki+urFZsQTt9xyTJGM4NeffynVv32ky/srg8PgXsaZgkE99w1ECJWPgQ4vn
gnrHxv1P/UjQQFligNUfjq6C+tNCV1I4uLEhAKLe/Ek3Z2mb+sZ1PcJCmffPOYIKHMBfm0+qHVAZ
QV2f72VFQIxMb5hI6FUMpG0XeBRuKUg558ncU0wXkabFMb4qLOsZ57SJZvosy4f05tlU3BYRJC4O
JDXQBN/fJ6zGF3QOho7olDnwy7xoyfieIJbznfJOTbSQkA5MrmhZ7EXdBfEPiK7N7xZ9WAzRzGg9
dwNFH4ZD1xVEHCgF7npSzz8ioNKtSbk379mSTUb9+TsEzQtShqpwwZwDAvEBXsbYpcWulYE5OjUj
PxjDUT2gJQS2b/zLNhP6aCOFJe6cyMAWB12g8hRQpFCOoNLlMYxaKyGnPuYLeQxJ++C0Nzu+sf6F
YWqZDkEJKFWSBXz/3E9CjMrDsd9MPaS6CYS+xft9mtH2MRjAdZfKCy0prveGrPNKP2w16aqkv2T9
B7A5/r2sYaBgBRvg0BMrwLrodQVPobmy8kujWEQcChBIXm6g1I3ndiSwzdm+94LbjeONWTW5YWO6
BS51acX2uS317ffIWjFvJVHbLwJdoXXy1wO5cWRl+aOrz/+JUEUFQQ8Icfu0sxp9nbpvakQcMmG0
IRtuTliw6pHqUIEmyThOtj9FgRWfE4PJ9DuUxiqpTtTqoeiK0xOxW2eoTtXH9I4WZ7y9+3VfOgju
UjYoJ3SSB7Dh24qDXO3FMSsPUVDKA0O6bXwgg7Yim4jNeoZpvT4sf03z/YwjeOA998PRXkuWGfLF
KFxXrHhT50PuGlXyjAspNJPP+P6fdEKCLQ8Zqzhuyotv7PRhZYXvMFtHjbEO6+R1nxCSeqU0LSCI
Wpu3eUhzwt0psH9cIp7ylbzhXHn0kcAvRZq78SNupxEycSC1JpHQO5uBGvM1D2kLMS14nUPpQV51
nPBlC//K+fFM7WiA6YUbnyNybAWxwLMtc0RkF3Oy5t0t8xK3lgVymHiBYFJ/rBmwbQtBmOcCYyp5
P5AUabl+rzoBSZZEDp+pGJ7oJ2nsgGaFg4RA2klkzdJBJQpa9yVtRERizfMgIcsudLSxKvY5Xf+l
oTq9DXpfG87Oc14S/1Miri3YdWlFjO12hHvzsPWJw7+gjLeg7a2isTL7/MTvwOeN4REQEJODSSgR
EUfJW2rgEE9hINZgI6+JU/4T4zaxNjFrn0wxuSoVC2Cmue8r/azzoCFFOqzdN7c10PYqd9FFlM+p
aGPRmBEqWU61wHFYm3yb2EQ1mQAppHI9kN6J+yBtTF/aN0FggcWT1l71Js1y/VKiYwGEbk0F1LMH
zp6KSB7c6HGYo5EpkhFnnHcHzV9Dn3NnTl4GR5+hEB0XzK+0QvaLl8It4ZrSzhhJSO6WBMWNWIaw
g1q2ZbWN57XoDCREXTIpNAtwz6A5C4hgy9c3gWNYmeAYHtD/d7ysknrYhtsWmG5yJnvHV6IOpYEc
Z5/E1z3gsj5Y04MwI90kiSee2xJgtVgEe/3f+SNmtrBk07u2PPsOgehX6f58fQhMHrm21QaqzM4+
UShsUTWcHn2e3B3nFt3hBftWyEWqEmVCgPx3G4juvSUXXGeim+Y2pgvn6oJxoF0zVnFhFFgOhi5c
VK4iDwVH+Iu0XH3NyNaP/+hUWC/FXogdEEdrv57gw6cxgwlufess/0DUsMUW4Uc7ggvRRDnGF8mG
FAenlpEjVfXlMoPA1M/eXt2dAOC42lVaFGb1/GdPJmVXlF57cNEgFA8uC2E0I6DjmhFNd+gH7lQk
uInWu6HjY1yqguV8+mzvyZEeiXsj8BjGaSflKC3SBSKn6TRPt26le3JAfzehg4gQbeWyCtNtojsg
cD04PBUWo5D3r+JQzrXfreof7srJHdLTyNM+lazxCHuZHnWrMHmq7qxfDoEOJwIDJFBpCJWtssjG
iPdHg1qV3buMvG7P7zJhMiSYPttkviogwo6r3cMBw6Z844fTTEp1lo/4+LnFV55NbpJIQ1R0RFUL
gl0K6/hsmqf5Udc4LqLGPM+RSqHX31skUYMzfb9o0uNwWYiiiIwmN1z0Wbtzs98lQSO9Auo6d9wb
wqMEaJO3ONhWcRovehS6kLj3j3mGPh9x0SEDwSVkMamlj+JwFKy13EMB09RXSUT7sGuLJpmVHZ7J
bo1koj1qazQZv7sxxSofYbm2Q17yCB97ZA+fR1S0UI5ZwEqQPQjtYRRVilGz/2JttZ/i53D/+f8N
XzGTyiZ8GBtZMeMfiHFidRzHrb5tmNnVuHQvmG20qxd5xe5bQI3H57cb1aLOPYI20wvGIVqos/rd
jOx8SZQDT8yUnQJC497KQ+NvSBFt7ZT5P6vhI5I2AYpAYw0Sn89uRqjihyt8vlXy7SJM+wWbJqzK
suuXA03wrKpqJsB+EzI9FZVkaDhS9sCMXa5SjS9yCNazS9xVVTW2fDEpNE87/S+ebgR3vysj6DVk
vQP3mbFDPUtd2SMAXfvG8/OMiEv/Jk3dGN0SZS0ElONQ/WDecNra7/LX+A/+pc2UyKedM1GWzdBl
mVOB20zeU4eFcTLjNSHM7rqKAcdHnl0i34nY1Wo2ltOEcfJWbOhJI1aP/LVSdHqFyKasewJBIA5Q
3bl81r7ACFsvG/k3GYJjTVfpSkBXb3kMuOxDOXz9XqX3HgeO+GcVEWPgfy4SE1sh0PkA+nEH9Pk8
3YAIAf0nAXqHVO+8n4SAA+2yCvfW1wq2H34hW5etaeSeJgi/Y1lyix1NXjRXZYUF3q2UuyKkHIb9
tvVqUwxlFml5VvB0/zqiN5HFsC0uIic/2wSvv0gZsoHHYCPMScJkAnfz7kX8TnxnXba+Ai/1TYqz
w9/MzvWpXTJihzVJOtiGdx0t/mXee0/kmCIZ7kualQXcxgLD2dLI8EtGYo7pkHsJKdL94taBap9A
SId3OJ9OTV7DFbB6y6NQsYo3f3iUHC3f0k04BSLQddl+LbjD6qHRbNcTXbjJK5DYDSHPqY5wpz6K
8D4JR0wMlFgyU9C/XJLLVn5k2a9R+3PlVnT5MxOlJ6HX834gtErWlzQjm9WMWvvuO1OsSzg0OsQt
Xf/XDTY8YFBdy4T9zwYfmZycykfxcT+1j3OhcJktO9o8E+L1liFqV/w0rI1e1gDkXk72yC1fMJEl
URcGV6X7BAqNC/Vc79QdHv13aRsk0OXHgr/TEplPsM4YwJb+MLrbcWhig23VuMrPIEDXr3tfVIts
aEEBRTjRlpPv4ZhsJNLFOjhz1soMEq3+gaRYb4CCMu5Apj6ifEOAopKJD9crDVeUsJ+e3AscvVzR
vlMgKDFxGenn9gbp2G9I/HAI4t2OafnIQrrDJlTIQhftGBmpV4OvvuoBS8QrclhPFBVhfStlyKzM
YXZEkGrWt0uXMZTN2CBy6sVs0ZoO5tRupMLQ8+0Zmw788GKs4XsA8FldzrOFiQY/7Kz1NEJDzZmZ
eh5QxH2qXUh25mR8NCWuU5IKr9j+8gEEmJD5nd4CQk7y+r56fPPS8kTKOJCmX1e/XTRexVu6VQWD
3ss33pn9qD4hUhSn/F0nCSeU4aQLyU2TJapZBiBRZs+W8xM+5S//v3Ldl0rpB5uNReUqJZbAdQpu
5f+zia5qWC3FsxLI+f/a897YvXyyy1Bls+KxihaYDo6Q2YJtFfzVWZ2F37qLiBXmqU2HAVxc3FmZ
SV8fx5FsD/PDZoYgkt7J8AuP1YULD1CsiZpvhpuz3uSkz/vtBhfWnh9wE+H5YiqStO7SyOGTp9d5
RXDLV3rCYWWKPbPkeONHLmxurwLcTHBUA9dc/doBLYV4pPIKjtSPoCFBffnbCwSwBx1iDj4EVmEu
H/MeMMf/hgsJFqLaHS3xxn6HfOJUfRqfagXhO4dgijH7hQbUEj/HWZ7NOW/9YzI3xUOhmwVhvuKS
4lYAvLnjBXwhwfHJI5vFB9EdUL73DjUvNsbNeYFdEJMFJhRi/5dNNKS4pWfSSoAXFswyxvuFVs9O
4AYldrz3F7EajlWA4G4dIh1UaiUqhmmWFPX0ori3E0QJ9+otnNAkPlkq3lBEzxo+RiyoskwP0xYR
4YHEXVrJDIe1OFDYgqC6vEOwGU24fkr5tnQba7JSOOVXG3coyDWFpMy+RO4nY5eyHg6W0F65J53D
8/SDGytzawx9di+NeQamM1aNd/9c04qvMe0QTOG7Umm2RWPW19iMHla3/QUp/tgQgTEG2G38124K
tE3RThsAEVliStPH3g/qEDyql3Sdh7qZYhUq5tKEzyTFWtgZUpG1CRp7ee0eKpEbjaua66OgofsD
XtKIWV6HunPNT7j8/+W0ZNyY7OaTn/F6OPYQSrDnBZ8FXpZOSRFpTpMOCVwscWg3rhpf+HxzzspR
4q/QNlaHGjuv3Dd+wcNdOkVX4fKG9XmvZsKve3W+iz0uwKrlOq7iqMvo/fsEN5ce5cHYomWwWotS
ScPhiy6bYVSRLQx7DQazXrMWg4KlG1Ql+32AeRiX2HM0Enfj7W+lStSjMKjHw3xV2qrA2XhsAj+i
CHEmjcThx9Sr/Is9Aq654WZeLACn5iOmQBx8Z7YeOdfcCQUj87u34soV7FoibLoSqdvYYai4P29I
6pGgudvvEZsRcHdbOyK+gDJHTUT2Y1mV1hs6xSGchM3Mqk3Iwz+WBhpBb3QElvWbddd/syUr3mJd
HrD7jKj7j0RMgN2P5490JIjUk+t4rRFudwNIj3VNLKCO8TwiAacPCwGWoSa+2wKaxF27hWbaIxic
uXvkYM19tY6zR5abbLc+zVy+IXOxO1QS3sU9qCsTLy8zp4hFStqV7/Eqsp8Mysv0Hxd8ddwNPAIK
JwZHqZTitcC2H5Cx71RHqo2Xfl9Me+ueW0+XFKayfSNhb57qLSLj2nzsphUQm2M1O3oZjachjfji
1oNjNAp58jergzyUEPfy+rf1RwlxU3ZoM9AN2gcO3gno5DQSNTmnKUr61jdojXfhNYMF4cDq6PzS
PIc5a7LCqQy1TBWDq+hLevPrZNdAvr6A2vhlL1vOmji8ENDIRcik7RS5eOpgalNSUs2tPDxC8XUI
UzYTZZGKtNesp3qOn3N74ZE+nid6d13x/wK5aW8xZNonBS6+BlSO6E5mq56nuljoRtlRk2yAJxEh
RbAH628P9+XcyF5JI97vow+OUCorvHDeTtOqRSk+nglG4BBa1ezSpprSvXFoCWfKpx4E5Atxo+2E
QRP6HvWAm/g7znzRb/mF/E84h7QWZ7GLNW3p50rM25/QfqzVHYxiCSrfEEAQb2SARRg0mBUnXI1O
jgSkhrhGDH5eN6FYLkCtl4O8Tj09/EssRPd98Tl5PX2JYq8FcoEQIRvWYTmTBMQdKEdNX9R+hQFN
Hdvyra7t2Fx23S2Ac7yi+JRfImBTCP/VRSkURsTky7LiINViqt1KSLBW1KsVmyP9p+Wie0uTLD61
J0zVEOl6r72bIfhKUjBbG5qRRhKh9MJFVFpJHKDxDuP8JAP1be72FJMOIeOMSeXTHCx1tpNOnklH
UlaLLXxh2JQEqy6rpw5fDGI/uIvU46gFmBCuITK1fhlYnwdRTEM02xTyMJe00i568sMUDXU1YlHu
oVlA9Mj8oMQPotESJOK9nxOo35VrJAFgcPJPGQcjxsTBAnC9wxz6XiRNj1rBkkstyWncDLLNUJd+
/dYm5aYzp8TWKOTEmOm4LPZck4Q6MapfmcF/pKaqEdE+wV72N2AlOIbM124SFSQ6afmAKciRj02h
ODvwvgV3vRbpbmzQ/FPV+KjHcLKpx+z6BCwEyf0/ijCXY0w7g4yeY+IyUvwKIkUgMCxgIY9peYV3
X8eXlGtU6bCIorTxgvHZeQghJNBto29HRGI4ErAeMvF7UXj/chpCZLMwQQyLHFgaNfAvF+O6AsKe
IYlF4hhGdKlq1gMFdcYX51+5uRy5u2/AgY1PnaW7wZOVyoaDOLKiel8h5wX3z9NDpSYj16jY9a8n
InDdYfOexR/MJNrWay+X3aGE61ve19+Giwq0pvQ4JlFs9F/CzWB/rS6ATGQ5/zYG2q7wD0wCNAic
Ddh/4brq7oRXvFUS/Rx6B9wFMGidmxTLZZeAte94apSL9hfpY439z5L8C2n8jXPROolhxnID2z0Z
NQIUq+Gk92AXmMlFfuPNP6m0PkPx1+CUrWlsqEF5vdpzCP8KQ8TnLl0Fgi55zUmEur/mF/mwBtiQ
bxwHgO2ueZBdAaJDyAHvkcjBX6F/hfRfMPFtOT+NQsRvrO3LKL8pI4VD++iYygMerVj1Jo/3YzvM
LjUdbF6iJkQvAbewiKuIk0T0BeFGukanbilF1wHF3ZLUSRhF5YxBNj0P8Xa5Fsun13L58aGFTszP
crqER47yNTELSIBtfab8/kwfc1H50tg9p6+3QpcJG0ZDfbRT1D/YUKAyuhkvoO/EutZU8o1RdtF+
mTov4+xGNC1fLAtnqpti/ne9Td9q3GKqjEw1GKUXCjcJrxeeh1pAM6+VgpiA2XO3rVfQABJEo1mY
QQ6+MZsEyondbAdiN4pIJGLa76tivFjpG1Wx2Rdw2+q9+s9CmzMtnYU3+axrIzqmjpD4cqJ3mwDx
ja6AWqKJ+zd1iupLRIr0ePi03OLDEJm5ruD8lWlTI8duwO3DWYJ9Kc+yofIBj7xOwA83e4AgbgXk
EIuGMnWb2T33ST3yGaxfoy0g+5ub3RF/Its8i4c38rhSDr2S2AHzVbDpuN9g7yBUKmF7fTRh2nrZ
olRt3RGUIAPt4NOJFMVUUY3/3brRerw2/qKyUHMjdaETKdl9F17t/XK41FVQD7NacYbpC9lpQPGr
2f2UX8w6adFgNjJYQAJ5oMDiDcJ9qzQftPZr6mHAXsBJVYYYKOUZeF8i9ex/ixbcRcQ+c05pWycE
VNB1AQv5fzOw8YKQCL83ha6EsqtncfPMu/XBghbGPY7WOsqeDIu4RI+Ab05LlJkdPYoGIUANPjKR
7TZIfcE/0SZIOGQ27QNR0u/Pu3huTXIaBULR0beivKk/0kDt/l3NkF9QqRiZkE2ndOU7pW+gNtwx
LNrevjWoYs6RHUP1H3RnND/UnS9+7tBwaGWezXC4oOOsAvuPBySVSxfl3LoFRNaTjWFG6Asno6xJ
mNGh7O9wY+5agJxqLJ22mgbel/pXk51NdDf63AIPf6aPL3NA7pFs7D3l7vSkkaZRTs36k4tSwfiJ
nWVBeXqq9WkHCSwreJWdL/l3+c97z13J2FoCgOwyeU44lzeLEJVaCuUkN2Y7tk/QZB+FtJcrtcdw
cSktaPmijxyt3jc8SVqhzt3xqRuof0zRWCLZWoEUE7nNXedgqKpxj39rSVhUOXeGY5+LTxSnumqy
jqk6YfjfYxxGxxYJ0c+UsIVmCBKSi1egb8JL4RjzMH8XQpots2+sfuzfKVNHLoMEzhb1XoJ6KPj1
hKuy4uKKdf/cEmL3LQHPQ7dL1hBkagRGzaDkxPtPQCw0U/Ht6IlBaANKRwdet0K1o8AipPiyG2Ol
z3HL9TPjdNt0E/AJg6ZYlip8r0r+fbhcJYA5S110MEm8B2Xt/e9Jslbxg+S8pFR0Av806IzTk1p1
5MCjNldOEMuV1ZSpM8lTN7BnEXGHsBHSuxAU6tY6BRfULaIMTPpUUk0m3QtYiEP/LoW5OxBvdnV0
b/azBWnQYHtssPucZcMw12pBqlzPJ1UJUY0UwpQHGFhRhAkLcvw1v+D/W8bC7noriLcvbd+2Qv1G
penrhzjaAQDGk00yp6A0sMmLmSsSlRi5V4ipKXa4YxnJ5b1h/UhTOiGCKMIfHhLEYawoh7ol3W9O
s6q+GiUtArbubVtOcg6dscidVY7mThMW/at7w2ih693kmiNySS69+J58s+P3VzQFvT2/vecwmoop
4KYmutAwPFob8noj7adqSVPnt8RMBYM1MCpBzv+U1heXjUqauzQ4d8rzPQDjMVmvonIxGSx2MDGk
vFjH18IYN1CH4RwS04DC6cS80FSODM/wjRexfrDDUAnJ9OoVfmMzacvmzXPN/KGIwHM7HY0fgFtq
Eg3oTlXKE75wdCLmCCdaiqEkNaFpyu2LkkaELEArXQqurLJxsDzN5kbRC01r2fJRMRjtospwP0bh
a3YK9ryX0dKH6zmIQHrYtG0nlqAc6GGuLBq3GsRdYgivvxo3lPhUa1rHhMnCJHa5J1zms1QcnvUS
n1mWQEuerK+hBXusj8p0firePWrmtwuhIQI2RmQ7JOBvpnnEG5NUdwRrChnQfo+fvh9FVDeimVxx
M7987OV4Vc/y2c7Sdn91LcFx62TMzDonu3LoxRSQFpZ5MXszjSX0NWVbjwh7qQJHC/PNDKFu7B1a
d6y3Ml7cN7Dpk/c/LX8oO0mqOSsBICF3FN5oVVGCsipVXwZVxvqlwG33uu5WR+p5oYvsVsXW8idx
maWFvjlXB9CllVsUOWq//6ZUshghWizAi9AtB26Q17Ql57h8J0B1RDibhs1CgJPTtedTtdJZrUWO
Zmtj0sUtgmPg2uyCwNr0TSZLSpCuZzOI6QnNaug/R1HaG+Qnd8f2tAPwuBohf5NuiumKBl3k/Kf4
vh0SlBHVl6G5PJBCYaZaAD7Bzq+paFpliU4aI+p1Mrv/EnFbDNMB5xI/zHhUHcm+9AwNcxQx4lRH
L8NzNCGuS1Vbq8gcGrtgny+6eOLINRczzG4x9OaK7v/FPS1Fw0nS4I6C5n7ynKXX4+mHQRcS+Xs+
ItBr/fkzBSfR39fZfB3G1yspCmRV9jiAaC4koQsiovy6XZfBRTnwVTLLmNbbMJ1gKzleTmTB1EyH
cB/31szg2Qw5cr2aWYtFmP3LEExOFWGR8blxuN4WuJrQ0aE95Mn2UTwIsAE1wwD7HfhGdC1haO28
28Jm6aKWnmzTvYMvjm1aJ/zLebE/RvLIuX3dLCcCWQMWqozyjhh+hyqaw++EOe/nfA7JnRGH44wI
dB1oIFl4sF4WJxs6e+rTBOC40leDpX6ZW1YLdOg7nLAfCMcrhEblqysJMDvMWQ6KNaywSsgLGzAd
EEKL3ObvpCuz1PAgTzIvGNLXPNuvuM4O3hH+VKCF1I1x7Y4fQTM6L5gWO7tX0oU8GQ+xxZ8drH2s
ls/6oaXqeF8dkdfHHUiTnyLUt8ToKtpaMVEbdx7skBpMpGgKB13fWHmRIjHHCPqbu5X0CcNdQIXx
CxEBWVN5+csv1nPhc4Yc1p/yljLn+zd0ld8Yvhjk+e4FYAMEr3sbVGjlXiZRMaO2fRQ52FZdmAIA
p7Ol6IzHRqypMcxN0dxwXxZa4CmocupmoNQHSyJt1eSOhULX63Vac4+xVvZra/dHAYu+8KJDQjHQ
T1pCdTFcZnYt4B+gGzGXJeHb6IeZFU93CC73vgdEEsUX/YpwQoPp1SLiRU1rDDXdJ/EV8frTp5L0
L0ql9Rd+wb3pyBhaWdmwWElmlhtmcN9AD1uK/PT4SodQbe6SEvvjvK6mOmjJ1WzTbU8JL4GvfUfb
unsTv7s5DjjSQZZCvJ0H6ndQNJ90xoZ3B9OnIhfqAEfdaDzdhb6xc5DYC5EXamKO4cf+Cw4scU0c
f2Uh+weQNKp2sUOkNQQB/ob/UXEJR0S0vPGAcyOUpywipyUAv/etzwvu+NZftaXgcNnollJhfj2j
PrDRrzMzWfL6gRs7++XZk/MFnyV5t8W9hKouL92eTvrbCLw1SuR2dgNmu3WHe8eRSK3ml0YnWorJ
e5uoh4pmnIPJGfv9ThU+s0HsNbinlonr8VTd8yyf/rcpiQZq2lTdxUENbBVTJjiOFKPyXQTsZ1uV
1sVe7MIqktRcuhN6qhqpLk7CPIwUY+svO6t9TPSE1r8hMD3qC9vhqeKSIP98zWlN7FGksg3gZXO9
P2xkdUt1uUoH0JPxfMPlm8ijU4X7bAsvSvG+gXycCmXX91Y8Lq4mAZjC9lNeXLms/G9UAc0Yfivn
vgdRamisV643iEEoDBweCe3Onr+u+aGEDtGUB9D706YDJ8s6Gwa5F9G3+t2NADJaBBQyrs3anWrB
67STJtei7UMXua26eAcjb4c5Zsy8ZEnv7AIeaWm5u+mpWABJ/zZEo22tzjlOWFhfP1sFDzoL8JAj
lzsWr1F/T3dZU46nJvfq8MqHoE86nLk20OqYliTLnwN+KQvF+LoNEws3RN2lx/CGtRFh2wP1XIXX
xR3nl7paOS9Xfs30JEPRX1WN+avrzoeIs2yLfYYTUqrVAr60HXHo9RI4YniaEwQojuI56w6TEUAT
6H7g6l/701Mn77R2T1eK+g2WemHHc+Kvz3BrePF/4JsmSrUkVjmTzldYtERLTJszmdnPxyNLhT75
67UJ+sEoOV+skFZrAHDHhHkjYaewX+fAE7KqLZo4hp4um+HqZKknNy4BS0AKHyVZZBBIGOB0woEp
NJMFU+3FT4wmfC42EEWguLXt3Wla0FvW7+RpS3CeuXbOnW0jTvvJuYNZEOSB/Px+f/MCWmWbi11l
k4ZjQ8GbVEkL+rSmTLLnWJEKKy91czEfWUlo8SfPSA20HZJsg0C9NCT2SORbxN4qKvYjkdzSTJ/c
nvvlXwxmTV9UP6NoHPQfl7iSXB3jV9zs+kH9qLx5f/6aFFYv1gpmtjHdMULNmhXXpgBYdbuEsOo2
Q1v9Ay5PYbBVmgL2DR32R16TDrUTk8qjT7EX8Nt6pCYW9Gl1im1XeF2Xy3dplbW9VAOPXITy0JBY
BtFSW/dZuFkEahcWrqJFRXtbn3g2gZAEqKO8v4iQmzBml22SLhnTtS188jYbb9bBAwJ9MTNrwsIR
Uth80Wuhsqb8z3ranVySb30HoTWSaIFtKlT1V9KxGBGGqRZzRg1URi0DeIWg0EdGnTOPdZJ5zf1i
YPkSq+YZpFcl5ZEm7RoChvLb6S4cNLMsqlWd0t9ro1rsnVnYJHV0c88Qel8JBioMogigXGHHllEO
Ho88K5G+KemaTJ9HgC5yk31WfayCHhm2kHRq8om4uQ8b0NqocfAiREoOGcd0uSl99fouF6f+dsPt
1jswRQBfekRJ2RfZ3nMnEUaH/V4cL++tASBSOyspuc2eVYADavA6tyi02lPYzMkFs92tG2mYs9C0
/5KB3+4bj4neyFjGitQmhbmVrYRZUaEdiRlei6gdD28U93m1JXCf1xU4qhY+Ut8Qgxrm0OCJ+wHj
fpwzVzpJ15DWUqEPraivuj/nrbuwXwXhI0J+PWy6dXIkl/EPhUQQclXKXvlggK/J3ZG0+t+mtdQZ
6v+ACUIM5gzs/eySAse12x1E+Gx1nTD4kmLR5seXnZKlFrHACnRGPZDbEvDQss/aOMt+atmszmAJ
7IYL1j6Rs8xVg9x1RRNvgqVKXptmmJhUCAYpGPRCQw11LMOVdTnahe/0NC1C6V98R9bONLjA8INr
mJ/J8VkRaM+e/VePnfiWjYoqa/RzTGnrD7DP9zcgaKGObIyCR65aDLZC3a9iU+V2hUAdPpyP5oFM
qXjJ1ZDiCda0OaP3nHT39zK3P5mLtimM8+QzRHA/T5YtTdZCZGVIeo+6FhY6P3JMiSKg/4sQ6U+m
ZpUGos4VkJ6YjR3QFRMhPD973RVwtuPyYj+D1gvA4xklcB9R/VOS3ry50FIjD8AwG3sQI8j83ZAs
5R2SEhBc+YMnsnLxSfRW4cu+BOGwCCH5+fFrER8xGc7H7VhZd+uFH3DQXxcKoJYXY9p4C1mQOURI
jJz9MWLE9gsedtROU+alpl1qevTOSYLHnOCaz/uyZ18CECURFgWgWGbUy/4K2zZBMtZR/ch09vGd
44s/an7zV3lyoA5TIEL1GcXtbk6MKuym1B8DfuKuxZidfaIH6a7HSwrGZeO6eYhNZX0ZzvNmF7k1
r3z0QrZhahEObjPSLmKx9iMMDbLSevCBhHfrDQ8e4Oejfdn4pXk3Opm5hKpzL/iVyngCVNEG2eEL
k8YPAYqqigS1GEudJbiIvbgxkrI99jZO9Q6dPBq2GS1dDbcjD5pS3gvjhIZAhPvIV36z9rVwtWCr
ODgInowBrIAGSuRMuaxTtJWsLO84eEYNWSNrfFb711NQeZaSb6eqGHWoB5yLIiCpoUIch14WJc6e
JNGHS9HpBJMsv1ugY65EJucZGI/nMfBLQ1trmkBhpz6fyblT6n0QlMP84ULB9+lqOFGlUtiR9LIG
6k5kfd4hNhb4xeywtip1MSD2+Yra6HNDvjoGjn0BWI/9uzDOEEN3+fZbMLMBPn2BA5fEAtxmSgfG
2NCDksiau0y5hFx3TM8zw6+2D2vNXrIyc2BArNQ+tyAcpee/ZwZzOSi/Y0nGNtl3ZecWAAZIasDG
cgaesZJyBYgWzkv0cPsls41fKgEb6UIIGaH53fcS6bHWgqCboezWxTiKJ3T7uskFTE3YibKr/yKe
fRpnFkZSOX7CxeW3VTbOQUAQS+8an3cLlIESwhV9n5jIHkszVDqsOZDT5H1rR7V0h1hz9+3/y8US
6JhlzpOgQInQjkse14e8VUemXWYBkajA2zsargVlyvx3JqS2bRzczDXIZjo/94OUvieHy1frbbH7
OI83NxLCj5QqjXdbdGvaJ4KyY0Mcse0jZY9D9OFea4SQAA4jVOFvDEsabVpJn33J0NvcGAMxwRsc
wYWcYjevfPIAGNB3jeTuWwRDYKSu7AHb75Wm+3EhRoZAjNhTVyYxmluhw4Ice43jNAYjyVslNL0b
wqtlVhy0eOgfd2HWOW3T9q3SP6RDY+CRYHX10ZjREtArDOI4lOFuobedBFrsuoI4yzsMa8Vei4c9
i0bE5zObuMt714j6TOJBZ04l9R7F+XrF3vTsioDOhkLt8HMv7/LKDTOBchtznuV/O3J6ByoSnZJK
KY8mhAxZTI8aOkMa/7Lo3+3FbmPYeovJuws+/Y8I04Ckr2wDC1I31JNCGc+DEkZbbZFx90SV2ICe
ckNUrtAwS9Cd2jGPZQP2zbxslp7lb1da3PSmqxXHYLveONC2HYDEEnob+rwwZwWf8L5Cn+6yzNJ8
FfiyHNaF0N+J5waUlk28qB4FwJ7xReu0p9bVMWby2JeB0AKnFHjfB6uwlgyjrwMX/cX1zyCpIMNN
i9wA6UBrAkOG+DSXkpc+B2e4J5KYzd0UIjNWNYRIX1Khutu48zPNHvu9aQ+8MFV/XXELyoQHDCea
+qE5+MYM14YazUJr0887TU7Ke6zpaWg8igwibQ3z9neINBRpE1C9iUXpOyqKjW8jZpWX2I+3rxmt
A46DCvmffA/xpMqXPlYeRpwR1iYB6ybsHARHn3eTAdpkx94IocNzHjwhWqxkrTx3z3r3UrYNhEsa
tqGa2L45lRndsiuEvBOQRmX3iZ6gBATNn24QeUy0Eh6kX4kJ3cSbDKTEySrzwl1452k3ljARi73I
pxjEwCQlMq1eVQiHBm0MqebNRJDpMKR+2u3I8JEFJFCtDGT6+LoOHbVDW32kvzfdOTlLp2H/rfXN
ce0ROGrLfJH1OcssakoXXOS1aP5crk7/eeJ25ydi9pHSCpKG0RiFasDu8DY71HP2Ym9fc1pV6BQk
aDwgWmaZxlG/dNDNT+V/CQXkEYyLtzcoLbn492kRfx35j0qliPZjBI1iwhS/1GidJOWueUq03C1W
kzzr3StlRSsbXr3xvoLAzuLVkoBvhz1x0LI01s11988vFtDtN16ImWlkMKixu6/zmq11Z+Y7iUYp
zoZswvsIfJiGqpKkPy/j4nS4RF6XfyBGVtT/KJbqCrlSNcnMlGSlB4Al0PORN7oBVSQzn9KHNxhp
wiq8BeLK/bMZo0b/gqs6JytGryCKDVeFFkIAPfJt04GvtNgBy2fnMoDKvamOiu+QddvsHhfwbbWy
fxqYo6sQcSZ1Rrvo4M/+faO6vDWNR+cm9zmFSXTspq0+YUM6So4C9r64h9nI8SHSaNvdU9eSPlt4
EI6l28HOS7RMrPIhCO6nXiFRj3aClTNHm0iJF9RawmuXdDxEi55TtDtX+0CyCfLkOPQKp8P3UtCp
3Mx9H5+kXjG9eER2XpFB6tFH9AnbrJzIEqn0Ra2iv3MiLrIZFCEaVE/TYWow6SNMCRMq1KHUE98w
0iwFLuH1WYi1NDutVlWTlgeCBPhBoJfPRviO14bLZFDwqnrFPDaarN7bnEtzmFdpj/u7T9Y7caJb
TBCon03BtqGnFY19LVw/AzXTP+zmxxOxZ1ElQyBrsALvCuooxWrRuza4iJWRv3+u2h/X+aSv3Fzh
JLHdIRIkyrvz2cJxz58HPzoBgDrCGAmf/5BosMcHYdqvO5WACk3jdXcv829hGXwYUaNqxDKBgQhs
nGYTBb6uSOAsyMODZQHeQYKmn8O5vq+24ZTG0pt6saZQxI8JBPZWMcjklcC4gDYZA+BrvenkXkQ5
IlUxJ47V/eutW6JycFzmYjEVyrv8xXoqSCaOL1k6yZe9oqgSDwYP9YxcCdzccRbT+xCGLvXaXHER
qbZnFahj5q5pgUZWHOr93bYzhwHo7KWZ25Rjz9+omAbGHhB8c5h2+RlTN81ENpJSbkTP/qomkIu8
3iNAZwJI7V9j+Pkm2CTZJ7kDUzlOMuusWT0rxipGCKIcvAIG2JFbir973/ekUxHA8dW9sozlvgMU
dN7G6QKyOtzBMFNJ+sMZT4cqDsLcjO56854COy+iGMj+4TX02OSCoQ5e0iV7tMAgJwK+IX6KktZZ
d/KT7gZ+A9dHD6LLv0mr/RrhHOVT/Z1gz6NZbx+J43QKb1wjU8d+jFlseq91St9mpb9+IHyZgBZ1
ppTHxjjBFr5EKFEv0mktSHRNPtlHQaChzlSUz9VjQBh8i0g+VZfw4SX7c4W2377o6eAOCHUR2AlQ
hHmwRsCzE5zVVHLfs1KHOI9+UcJjoyfg73jE6h+G2TfNUGBpOluouC/1L8hTvQBjixsDAfjuMGad
l569lr45A6qzCoaGiD8SfTCrU592vFrfLZP5GQ62cTKxfrmD+3aM1isPtOnT8nO8XAt8yqNuiZ0v
buFnRYgQu54gogMmHHWzkv5DPD+3a22U8jZm1lHuw/eBFk7FRozwrnN+Piz9MENqEAK3V6eZpfqJ
Lp4pY1CSNS+h3Obws+PgKyAfKzDYMktmKib3gAuWdxr1krqmk86u9atuk9Sj21p0H3QNeeVQQ4Z/
Z+cZ+SU70SvRtiIkc4TlhU6jtRbDCAJ8gQ5rp8LcDBrPvU42JZeX7fXKWjfFEUVjpb6vS/5YU5dS
vOulItEGPgRdJLJK/2HkjH07DpIsXutlLSG/5FE/PvZ2/X7D+K427cyb0mBpaIA6d/3XFvgSpFS0
Gt0hB0AYSzPFTHr2e6eUxtNyJM+HT5vfSnAM2xK3fBfnq4JBjeu9sth2D1/qDT6NfmVgT/wrBDhX
ZTzLY4MihSxTkOcJ4IF0Gket8+adz0kRaZZCMByNbSxWa3D08o1BRNsLC0k+1d5JLNIV6RWnY0+Q
DvCryMMYu6ApudwNdX45AwSUfwUCiVz/ozRj8A+pAh22wpD9/+7/qrwjV9qLwWnuzwZkd1uLFEyd
8I8u/Wknakt0gwt5dNIwJcdMsw4s79dDqPlCULqlAr1Yw8fhzWszNnQnhX398pzY9hEo0r2Bki1/
HRlSTJ21oibaPoP/Ajje9KHsNFmx4j+TR4tLlEEmVoBrfPR6ZFodiWy11urq6hLpBmyv4YdvrnVY
TECIUPhMHrlYYSwpUZiJBTS8cO8yfBm6gjHyLZduic3yflEc0GRbruoXx87ECOGCqKPtHAADIsji
2gZI6MIuWjtzY0jBNrgq/9mOtfbTujLttYeGVNRQ4GeL13fyJW8uGXCb5Ok6rsy1N/MpC+uRmULx
bXIbTIV3tPQOKq3jSkdeo5/RvEKKQ46+B7MtNxLh6NdiyGqetGAQ9LyuEOM5BnDdj1OnXYV8rkhs
xE1cX4E3O4dggC9LSMkDvsOL0DdRgGAGFUHvaCZyhAfvcpJKERHvXvBUssqmKt8VJl+56fUjEs+z
tiK8FDSH+a3lUJ9IlmQZBHYQeq7aw2C3lIUaUEygnJCIa9Ki3RPs7ziXrn3aOxVAMIUyjNjMBjxa
CkfHUkUIX6QzmH8NQ5KlIhUwXY6hp3a516gb3q+XqrJqIQsseVR3i5e/yO1GPIOJ8y0JX4xlIyGu
MoLuB5hE6VaAuQwvPbR355Ks7xuEvuqt053kfjTmEGV+A4Ap8oF+H3SwGmlI1UqPv6SaUdCq1lxt
3lahaifh1eoTNjEFDBjDJsaSeLYpfSGQNA2sEllV6m8tvQ6IUmVdiXbsnEY9BSwVjZxeD85KNtqP
WQkOsaEhxJL9cUzHqM9Yl9QPauzMDAKoiIyE0FL1JpK4ZguvItQXEoVoR4KlxAIuT1uuJcvftHm7
w+r7GQt3ATeL+m4AD3uupLmqz/ZXOONAJQz/IP/K4Kabfb94pBA1Mm1pddMCKygz3MBNJ98YYvXq
FoiI91KfFfQoFRJCqiRqF54KSMp9CUL647MKAuHOEp/lmXfiR2Chz2JkvdZhYare3JaV0ImTKgus
r0Yhk/mlCGt+nR5c+7OCsfNaffA2Wg5+zn/ejFMCaBQ9HZzBAyo35w6NdL0rU6iYbPGK8nwleSNP
Qa0NYPriNsa4XiGbDaKHqIR6sen+enifTNsv+vKdhCzo3bHDTx+vDgAzT8veYc2AUgMeU9azx1Az
Wlpih+jJfJaxuj2ynHtbSpxgxFVx9C676QKq0fufmFAkJ53fcDZsYaRmQZMtrYCTupAMKYFwIoJu
6OlUcbIvZojusI84oWhGRnwWK3nC7ZjeY6W0DUNtRP+FS9Hgf3M5ui2SLrVcvUCHdeNjqL0FbeVE
+ONZFdmxXp8+KZnL/uWmHWAcM7RoSKnMh2Kf39tegzyF9BiGvuQEGgze4lUZKb77NVD2EkB1RSX2
wQuq/LnY5eEQYaqnval5gQ77ysh7kuRyUPAuNAMacuJLp+/6iPAlN2t7gy2nm0BiL5FwhH2Tks3+
hvSwdOIxd4Ce3QXO/zyhHMEsyRTOWbfNRXZbcrz9liIRsC7eQe7HI89hsReqVihcE7gNXFenexuK
DhpSBRb+8TzciT6/Zk3VRrxUWFUCcWSG1Eq3U+HPErTmXb/0Z/JTE67sVz5+lu20API1rO7nYSUB
NiQMCvJ/98UsoxgMb0PZTMMPgJ+vlqZy+GcodBuHJMK1f2jLmEAPxL+r7JzWrcdd1FiimDhSKIWe
+Zei7c02aiUkD4zwl4gM+X2KY5ob+43386iqn2WNbHSR8hXBTxOPfWjgVIOuY0enn6olJQ5Np8pJ
unC2Xm1e0it5IERoo/ZEsc4mNM1El7hkPnfnHFmkOHr7T2nSliAv/jOn46XvVWr3Tcnw9USwDI2P
g6r9xncLBNWSwaq4OIOnyy+dQNYVDZDGsYZeaAOEKkfQM5mHHPKActwrrKxnHcTdekK4KGDVI81W
yGAGFNOLvT4wfMNptBN+XXTPmgd/AJEG6iaIc6kF8tANwKfUvclr7QrtZglLQdD8M7Eq244TZyUn
7kXZV5Jdc6loY2utxxX9CNiUg8dd81hgzk5inew+W2MlQDZmr9A3t+R7do01ZVGli4ffAGa3a/2z
rvV5YbWztdjFky0xhkg23unVlzk5HaFIgj6BgSjgY10HWxz0oOFCRMZGTNoISMmkV44l4AglnAvR
nl3KoAXlZXeiiNVw+MMCa+6+uy29G6YcJIqL8x7OXUUSN3nIymaI879a20/NnHtqhWzebQ/SMV+u
edaNe9zU7VCzHDRr+8nc0OZ+fpLyVllqRv2D6ItPLWhTNzpy6Et0fx8+lFjA/+IXyNSb3swwb8zX
RYrtqaLUR5jgIUzbh6VHFxxPRnXOie7I+YCROk3cuSppHiRKaOLVSTx+x15oU1Pd2sOmKK5lcAcL
Vu2zkwYGYd1OS9SyDcxobNW0Zq4MvvjjaVuQJcWjW+VE1VPR3zLJS3Zp7vFHFMUo/TarTQzNDUhq
0a+NOSOuWXb1igMJ5L+rXmZh61icTvsrbIUwt/jiezdFDcX0Ft9ar9+Vy03bqN9pGgAXVMOXJy2/
eqXE24DcmxnKEhfAZirjE6N7D5R0YdeStn8ZENZ3/ir2nv8e1agsLLfQUi3uxGlFt3g+4/RuZVNt
3rfFJYK2oaK32t+s8OUxeciwn3qDHXUKbJacM+l1krTa+fIv6NWnh7OAi0E6UKlYm8eNkJfsaYX6
6nwapaQA4sXZV67igPPBcRp7YLatxe8DivILPzj15qO24XqsTO0hkTA6wBZ3PMDQprcDxtORuO1T
BGGBeJdFHzZUDrrF6CE/OHeI5uebmnulbLGZziJLo4UGKEGNyYWhqkO0eXb4dc5eCPjBC6qnUPTv
sweNA3b8h7Xyv5FPKVLobJp1sAjvqXMpxcuv9VmEXRgEURHwNGnN/5hEod4iakgsVnj8vL+5LhoM
Exk2msWflBw8a0OVxkxxG/WlSpoyXPbyIAESLw2pLe7g0Ufp/RLKnGL2cqcxSe2beYQG9Z6qlDrS
Dn7qUdmdpwmJEDuKVQA+E1dPYQTPsaNOfAIVVBaISLoYx/gL9GjYFaD5W1VEmG2oEtNbdPLpKv7+
SGmElj4dKJCohZCgdfI829BgdPKxCYcf5LMLJYLxF7pNSuQUoKvEIUoU5vaZsfFRTkusS4ozKs3v
srvmE80JmosOvFdaRy9q2xdOGUrHa1NJcZSy7Rb1ITuTLdwDtpVvCXBE72Lioxcvd9fKZboyg/d7
6tBvK+rXz6owNzao+YMTIEQ8o7RCvvU+0CkZzFypTodbkocKrD14RwPsOyeGAK9b2MWKGFNwgqrJ
Jvhubx30vIqzQovl3uu44W3HlvE/ENZi4RtlYizLSxFeN8lzGjX5gxYqdk2bvW2oKmmXyWkRToog
r5DC4a54PhLpCdhIS0UUVVZdp+EJBMQePtE083zlAx3pRUkPVVbVyCUKvxAAQD3i9DFxR8XykPZo
iHOvu3lvVzLKLXgPy4pItV31g9cGkG/CUc4d9JHakNLRL9fC53Mo7FWRuy4Lm+TY6hjIKUMh5azk
vppzivT9tvMgcWMkuqAIxDN5YPyKh6cFVHHXM1uKUTsVOVR5CRfsMJMZM8496RnekRHmPB63LO+k
C2Z2VYpbqiTzhWCQI2CxeFlE9ZwNwyVaAaj0ObPhU22QSnq4Gpw+ma+4ec38gLDF0CY229KQzy1S
F34QQ+7XpC2TfhiAI3kGw0NObq1kKIc2NY7Nsyejyt/L0teAINuMrWF30llsIPrm6vVw9bRGaRUd
Z4NF4Pp9Ec0BJQfw6u0XtftXfNeujtWUqPUN8SRiAVi7dZqy05SUZnBJX4ek/dw3i+3tNz/6ZARp
v3fLqXbbW4JoRIxN/JzC//V60cxysThVjjmV2T1/tmzNVX6/1VOcAyiD1g+rDtPCHmcdWVve78eL
YqC9DdqUiRll7cAdoOzVVlZUMPEXiJkw8HpClnixnjKRF7MIVjGtJ+Ay6SoE39T8w0GYzwfw8J6Z
5VbY3M3Ncv3cL5lVRt9C5IkwAoZdC68+K09O1UwzvS8RYK5wCk3Oqulsp/d9zGPaekbCdgJWLFSq
XfiCpgaIrNpjHwi1cak28Hl4/Vg3KEX3Xks/lwj8U++o2bKRL5TkJacKqilZEU21xzqsgmfSkZks
pK3znCSHWY0IGCub1duMuuloHwbjbPtY3HiJE+aUYmYkyZLp1EzAxSlNj3Ure5LQkrRlP6hviHo7
K5idwb4Eh5nMZ4ojEroYgwoCCRkxxVGpNH06W8/GciZ1I1IT/uvaMtbhfAoTor56dZORV9vTexpr
8Dxtp94MWKPASxxBrc2/MXXqH0Ds/frpKxmBvCCv5rt8FBbzeOmee64LPyPWlwt2HTL1paoEV65N
u02PQhcEGyPOASKvk0mcFEK8+fqJHgD4G9vXwb0KCHVilvRlRJMe5KJphD2YdvU/VBfFCcd7Xxvg
+2K2NGluwdUE2QndwGnYe+KenmWMBYjF4Js5tY7UOdi2zR4MfQhXfiN5CquoFJonZAGTT960kS2Q
hOgK9JGUTTxT9U6/t3TefngVu+InaYBWmaklDYtVXMulVD6IQokqn7X69wNIEuc5mytYsXBaYzoL
G1Ug7RXyJl3bz84O4tJXem+M/3DAesWEdBJTsyHcRovmC/MDb06ZDY0hfcxJEhl864pQJfp/8BhQ
7q/f2uiglI4fq0iAscQeV31Y5hdk8/d8xvNMKvKf55fEZi/2pCrNWOTOE+pO93hpASp5q5BJdHIh
33Wi9TmeuVwzRjy4ZrSag2y+Umv8CocfP8vZjGdfzrfv5z+9lgSQx/MgY28zN/Ile0GQJBVBBeCB
GC4t0DeYYT5gQWcNYhmXdaa34mydiUOUCMrxhcunA7A4cAqqPWQTFp200Oa0rqFe6hoOdfZPOnC3
a03oFazU/YHOPGLEFN4FVi3P7E/vwYd/1pLTQmPIwhkIdYFcMQ0LJhdQjxOBs3mX1o46KrL3URTT
BrBEXKQZEYTPjPWQYLG7ojHJqpmFElGFzr6wIInJdV3SvTU6xvj29uUmOdXYPL4XlDw4nrMnHS6i
7ZE2EvB+I8CMsiKRjCndoEwLLUbNZddQYnLVa0CuQkGQhYUHv5A41xysbhQTMbGQVyOZGwbSmGYf
Nb+vfaYwMn4jKryCQ5ciVi6XeBa0VLnrJYG5ZC9UclAssXsT6/4gexW4kjfy1xO7fiGc6HVhoaR7
xN+Y9KVC6Ug6x5DX+6NsBCKRzTt2k8fi95bPJ5+2GCdr4OaL27noVVOWx1Pr2t/ald7wPT14GMsV
8lEmc+PNNPJWWa/whNeFC3LOVrwa8iKyVwZ4bEeiXxeV4b0DLH+oZTg3MsEEuQsPCPJq5fOIjipy
dQDbPe4pMDYzIgqnfV+pI6MGbnQG1N55zE40/9fqaJ7it4z5ZXFfKKjKvxLD+B3z5egr/1R28WGh
zfaKKPn8jqUma3j4OHfcqQ4ud5QQTQtlpwO81uQyQ+Ffw0sYQiZKZfqjrN3Md4UUp/89AelxuuF/
987BLS0/k88GEd2e69L40vh6eeCRmJbTuL9bF83NfIzxNTrfgCEeLuiAVoKeihUEKkuihPyFLz/P
8Xpfrin3xtkynVppMsgOfumNfKLgM1NVC09e/oD7xpaU1NDb8iYgi9+6Izc9SfQL7a17olz9XkQh
IbMJJ2Qyp6MXE/3JYUiue/ykqwbs90HvpFWfwAK/+I55smgsFBrKigZ6r7Du5qBlmLKE5m8p75x6
SH3jv43pRIlLgf/Qi4c3gliCgG7acB4384FZcV/9TxzoGbLVU28UIIZ5In1EzywG8SFbK858AXMj
2+NqF70yt+eg0GQEw0NpdjZ7fPlfSFOVsl0hztug0FmXmsmvwii1D8kXtRc05WJt4OpaZ4buLvXb
ZLUW2COmkBWzUnXZr1DV4q/RLKlWzvhz9B8edlo8VHmU9SA25RJeVEGoDy+aaJg8FOThIegqhjOZ
fKOR/w52Nn+nHKRShjATe6AzDycWkUVjypuo6SBY76UDdCKSLsHnXwkpuaeq5FUqQFZVTpxRmIvj
bFRTr+Ya/461ZCV7n1PqJb63Rxhy5vgAKkckBtOZ6ovbX8Eu7OLBU4izxDcQTjxKu+FakbpspasD
cryv4zt9dwyabKB+pfj5095fxYlpSY25eefEMwKgK+4jvaDc3G4+vFrR6d8VxhDA/9GDiB0bu0Bu
qhi3XOc4a3ChxVm/ZwWMJxqsWfiQOOwb16EbWzF/iIBXaS/XZfmgCHNfVjRcEd7PjFubvo1CrXZJ
GEqkMSKR404R1XDAB+9vMmlO1zcmilXaI+iIljGfJvodsAZKD9v0btrq/aO4TI7MKNnLRwaodgB9
C1cC7CV2CCmPxKzt/QQr81L84TbGUH8bgXHFHDaLXJju390G1/AalvwmN1OmAmZEJI2Nbp8XgMZE
BpT1Awcx8SZ+B4EOhIKpt7Xihltc4Zzmrj3hupa1gX803DoGVcCOR8CmLlXtfqryUWrC5UCQ0u1J
Dyk5mYwpEi8t+pQJ+uPjkwUr2bAgzMVSS/NUqPsthlJEfRdTieOwBZ/gZP2lUJqzD7Ehmi7Y9pje
YkW9aSjGEH+YohgTelfc8bXZKqXLRk4zA1V0owf0oy7Oy6Vg92nfoUH948IUdI5erKvbQj1fIOf/
7QxDAW45/CYUGof1tcUDA5CG+N4c3yvOJdhsoxBIM1+zkwpkXFHDCVfuMimNmSAmtuZu/nNydziE
mHX30cImWviS0CDa4jyMb/IL96Y6uG56bpUdCvcRF4QVezpD8n7VLleuuMGPgoq8jJO81PJfkXBo
cJl2SHYBcfnPGKXJGYWKla2DvZsixLrujQP3kShr8oZHA16hEGX9j+mSzctPvmVOYz2z7+NJgI7U
WNvdiLk0x1st/MqOm0l3p9hLa6kaNrvkiXoWO/mo/K7kuWMuwdlAT1qOEQUNkaqarPWS+1Q/sN7S
MBodrI6fG0imB+fA3R6yQzi+tJmQcbWSwk83nXR5O6+UuXv9e+8VjKRZPfKo45ftacybGpbfajb8
1P4LsPdkYLK+Um7JzldtOWJlwJdhzKtaAGbVJYDZHfr+RCdvGTMfOLRsmcUAakIVsfalGaC989PW
mqB7gHSKqaXS9K4xDjBvqIf02oiKYscTKs0WGgYD0P3mS8TtxRwICxscMPqghVNaOt43LXpwnE3s
HaWvHijkiqETjc9AI8VwKYFFqdsSuLBbNm4GND4Q+rT81cZzc3Nf39SW3As293QF8yxTXxypXPhS
LfyZnxAeZ2qI7z5xIWT6gVEBEVgQ2T6UlpKUCckhV1WhHuij0WWg0NOALfpOjpAjRXaaNsT1wcKF
UZt0acDUOTQcalQ1Of12nWAbqOAyyhfy4lGHK6HtsZWiSLQuU9V5UbtfAo1jaNnguy55giVVzNex
reTtKZRnTz7kaARjQ5vhAbVKQbdo2n2TQ/Gj8/XUFdxS5rWmruMc+noIgPbNS8H8vyCpuc41dcYO
vRbYe/FMRqU8pZH7X+XsjJ+9923kB8qJp6qQj7ZtTE9MQzAPkwUDAyazfn9t6ymmozJui0ey2QMP
kDEAt5lAKaKjI3x/3Ta+vFgIYfqURKRAPKnSVbB9uFnG+Z5FUilNzbBhk2VkXs0XQsHPgDpiU1XL
K78Kg2YgYho6W3DVema3vqwOUdWUt+bl4LH7NqbwJQduAposlGG9aAKsf0AXSyQF/FVcaFeruxXI
Szv28/zI/4gqUklYCmP9GzBqo5y3O21jXTNu7n1NLFmoxBK/KMGoXK3a30dvdYLqILtW1eevMjCN
5I/WE2UFC3OGogl2/zP/hQ+LhlD3oYb7Y7WmUk2o3LBhFireHNHAy5mRsZp8ODkcq+bBqb3wjlir
3AJW3wcmqzlZT3Ja6zfHrr+k3sdWSPwEQIx0cpNiQ5+VpcoxQ3LjVAQpl6kDiw++KURAou8c1YX+
D5Z+tgpZmgXIgu8dV0DLQ246t0aaAU5wYlU5CEyBTXdAdpESkg7i5c1bronGuIrrtpJJ5XuGGzLZ
/0maHzL72/TaQWBhnOLsb46jX+XFfSf2bdzABA3fjmPAw75e4TONeDYmaaWq7bMOwoVlEw/7OEQp
4ltO+AAvAkMR1XHvjNnq+Pgk1XSlbK6UB8nNhGMu+cxq9j9DdLGxK9mzlfjzO8yPF9HQ8tKCEndi
zH4GHjXVb/QPqiVBRDwYy7+pHvsWsZ13amKK3j/s2utGQSKaXX7rIrOkTlRHkd73yaNBU4TcywPQ
Z+/E9IGwlue2gEr6NMeAGg/tSU3QhVcwDxlYI77w6T8fhaBhZKe2GVVJyJJ/xS3OoSgCuoTRm7MN
H4FarMCN2045slnBPThLeSQz3Nl1tQ+Y7GxWAmY7M7VGLvUFA3cN7Tb1LWsln+1S3SQDwyoRV3ht
iU4G0slts1nuT+fNHkTIVQsfRwIkcUm+wAmDaYd/Q7YMHdXDzihV7/5j3D3JJxutWvmA474wLkHO
pjL1UmmTvTdtk16+fj04M4lRSbn6gqYZCbVgHlKsy2lVPwG/nS9rwNAXhskm8c5TVOTzUJDaQpBE
iCpxXz2M4ANgjRe/eTbUEW92Dqj7etBXO4JpaYgIIP7d4bY/4uaZ2JFHlbXvefegQTc8WaoYkpMu
tYvUXDYQ6nOEKWq/87wokk6saWDRkqDZqrvGObCI5AGvFZpXOV7tQXW3dF+UEdqXFJ6ejHhB/gGw
Wit9MIns6GanVD2gaI8mOQqTSkD+piRybcX9aNOLWulU6EgIYl85BET9gs6arMoMvTzLyOv45GfX
pUMG0lepXuKVlmL95Pp6oaScMslUke0jV2NCo4SH+aTbCTVUASHKFQMOHrKCaxkhLr4E0vIfCbY7
/7OZu6FgRBDEKpgehY/3RZbvdSvuS+nNxl2Mk/pCpk6CMI/6iLqsnotUhVF1bhv2HZEr4GErt/g7
1UClutJBaRCy6ChhiPsqt5MMdgsDa3syZIamnZgdTPw57RLykhYsgTN+Po59mMRejmzpW0hNssPG
mcyK7xTAgoV34kB5M2nX9uwshhCCsSkxr9BLp3FGx1zClxEp9i5pxD3iX/knBRFe0usfhu1ZY0M2
gOfFlpTlctYheehBdcgiJDMAr1RXPH279XNxoYTPUgkMOPTGqJzIpYhiAJtKFViKIIhVMfTFZEeD
QQKZ8FyC7qa/z9nyrJ8ONjO9H9WXMr9Qz3vN++hrnVxTenS2S7pqz4xNdfooBmR+qJp/KNwF5YKc
tOlSXYwuVwYYT1SHgCmY9a+T8ej7IzqRcNrpgSI7DHkuO2a2f3Gd3L1vZFIQyQnIxhR5vuBuxwbJ
Cz1+SFPqUhbmci06yL4xLJss6r3pFkJK0cF1w1757ic3kcFLASwIdMs1O60VWqn1zyMJTUGhJqdk
a+94owgWeVhtnClXU7InjpcDrsbogvWKajTqegdsgBvfxU9fyqJbCbKqz9h8Jhz4fnk8VlbKOg9O
W+OZesPeCGpJ/m6jP/jHXm6JRHmR5u+njq/VK9BSWhtRyU0I1P3oBVedccPYtnFwiCyP8gIwijcl
evJOdNnjIfp1ySsUmLUHKeWsHjHVqvnSpIwZQl7ItiJqA/EYXuZgLxRWHFMdaQShu4zuSBc6WTOi
gcFxEhqr7+8Q3IHTT3IJdV5fXsuALOey9ta+qV12Gkh/yap7nIe0UJCiWRNjnQVyHKrSqfaOz2dj
DJVXxzh1Einqobc5x1MmwsEf6A1iqm7PsG9+oP1iIcgpiZQn4MLIH0cyzDDXipMgfnLU5s7pL3Ap
ggOWgih10eDA119ggVjh+HF6lO50GCJji1jtr3VRKL8IuDgIpWVspXHzSuyt73IxSoUztkRwSLpV
NkP/rKaTZ3zClsPvOkKG/ImBJyAjCjXU59WCPj3cVjrgIG0Q3lKw45L6pY7N6Kjwnaki04fn+ghs
qTGRZekBKXA6xTSPsp2Y5BZjPz3YWdVgLlyGJF211Y0Bafoig8JKf1c88VM4eeI5sk3krqKYjnvM
iHc0apKvKvr3S5ZRRgORerJf75yeGXaGLswhIQ1RBMyTxGg/14BCK0IDNjQTHBnRtTRcQA/OmoQi
3JBWFuy5rMmnyBEZ0rWSPpEHlCaUuuTBzuZB2m7kqPwtTQdROpR5TBcDHbVOL8v1ks4D3nnsodZF
frH65aQYaxzfbuFHAmRN3jDPxGT8shYF9rLo+6U3CUApr7BGik9ABDVb4zG4pyq1VcorfqblJFvy
lwYxRcsNAidJ7ilUicYUSv9h76Zq4iFAO0or+80W0wY61udHz17bBaGkdqjtHh8bQIhApJ56c1LV
hg16IW6Zb3Nt6q5Hgi6XHwzRAayGDxrhsMQdCCbqiTvjlMc2PFdFAeYaxIpJ14gtqhSh3FFJkJE2
WC0vm61VOlevq4jjI+n7bZ/8LULBbWu2vymBqqvmBUiv2al2in32e1sjcmJ0ywfncB0iPC1+AGCh
fJdfyKCBFKUoTaF416woOEYZbX+a8hfbmOI2aHNzUk8CTfHy6oqzujA8Ybx/FoonExmKE82AsFyb
OpBVDNo23BMTl2HhjDQECvKbRP2uEWGgeRakzJC0euAir7TOR3gCB3rU+ZFHGxAOPy+CThqza2w+
S0t3Qi8UhwZBvyq4BxJ7t6ZafrYcs9ZRS61TYijMSDorNe/9xZyrxGEY6R5edLoDbEmbZqkF+KTo
n+viN8MwdlcjQN9NNH1bdqJV7/1Jfawc6vA6AX5T0yE2vnue8BMC8PHHxaieV5xapm5f87C/92m7
j0bEEqHfoD0afwZLBPromPGOxwiEBmSPezVP3CbVEiVDrd2ltG2hsMmhfgxYwZSdc+Ek5V6DJgE0
VV3zXDQpbhi6f7ZegWbDQ6njI/pUOgPd0/ov2Cy7dubl4krPd9I10TK6bnS9YVv8gNOeb+cE/+39
6AaxT6fEHYAeYWGeGkJg0JdgZNuc2QEW9/DY99cKzDZsFpFW3CUYAgLW8En1J/jp1sP/nnF20x3i
pOpBMcR9cmprnTFGXMd1TN+zXGgj6nwtiKx0fF1t+cmNM+MaoZfVpM0epgLk55e1TNsuF9DdyPJG
0rLzBAVSnLzIDMiH/HdNllFlSrAsv0Gu/G/OkQfnSrZ+RbsrzLZKWfu4Saom3hoZDtOKPNbG8ur1
NmP4oH3/CyzjUTntI1nI5arIYPs3WrHxKB17BL3vGZRtt4P27Yq4xr1n4/e4UOAkQ+TXlFQsqfIA
2Ji4GN0FAIjBWSbRuNd6lz6dYvj6S7btnaCu1mfMGn4PTsLakQOIPpQ6ihw/x1K7WxeTM8aHiNzx
yk5RdWtWP9HZOcH7kIELE+YfvW4n8GmQDY924goFFjy3pbzxnXTuNMOhi7da9qUv4SCXGE4sJtA5
7DLYux1+8cvKLtjU1O8uJP5mxgeLPl/3L8sVDTieac9siTJWozCBUWzmXAhgG85q6uR+Qk+SW/up
txKjcLIhTIHkdho/jiv1CkWLXZ+YOZEmoZPGvWZQs9YS4vlaptA5XbYUrQkPbfSHQAjNXZI7VxAa
XoL8A0p9SAKhIGLv4q/Kd40T25F51wTZqZkCXGMmea0etS31m3Rag3+75JAw2e7IVj3poBHlEmIY
DpmyJms0xUVoQjlY+AwcaE0W9zbxFqnbde2lUReQjL6jeHdU50haATDACPoAh4EGymUkvIhDRTna
XhpHus4oUDyEq510+f2qHT7UOIMY9WH4ZarCiiBJfjHC7Rp7IWEM1a80jOsmvYZEygTZ5ALBMyAk
wk2Tgd4pOzh68cx/SgfI044VWtzyqLZ4K1rfeSEYoJerbTX8LaM9uJjXNDaoeJx13J/+5bYSkNuE
WgubXjvSljUZdell7Be2pom+79NJBZJ5MWUhcx4l2qKN9G2ngttsya899RjuvoQ4mznM3DxBLqdZ
8Sz6uFHqIonQOLkUR1DqQqAJf8a9bAKBgqxV0oOV+BZiCg3kzfo4PYcV3Sm3RE60GIBccEpbUBYf
sDLgA9N7EgR6icKPxs+Z6rJgcd66FivVzfubjdFRZhKETeSDMOAPJN+SDdyeZF1uhGK92buIjPW/
1uTEOJQ5kQUJyN315Hnmuuqbe3oOJPT5gsxjXq0LF24DFqQmgAhXlzlLMrfsMFTnL2RLn9TyY2y+
Pj2FcjAyzzzwbqPukJxtmlskQGhKqqWfkxGnSluJ37zBVyf4EiZjeiV5Tun20kon1Z5lLnTFj/86
dnqZ1nq8WNk0k+5VXIFhbNJ3bDfpUawHhhSMdVrozlSN+1qhy452OeC+dGr3XNj1WhCMy2J+gvnd
nzEBe+itmHksZWh3ADEyHN113Dxsmd//zS1lPpZNFV6xbqReZfg0htpgncw0KITfvaxvbmZDPHVV
OfJBHEB+94nlG5jMgpAvtN1J1vm3xE8/i4I6LcTcaTztWUBdMXbOX6njNwjCV0VXhj00CBvES0gT
Pt9jrLbl/3QbTmeGZeYxQGGwzv6VO0TVlLx8fmTYJPJ86aKFKAGn840/vwyXnnz8JsNG2zguIjXF
Ed9jIEuk59qoQ454ZQUltuNdovFVF4qswYOtOh6XTNMang7PIn+w9HX/dzpceZ0lB+jcE1PpyfQs
wpXK2HdjZfgjxQJTYSYjyfRjjqf6762ORTK5OqoaIeAQm2pAjyTYH7wRiLTfoJVdQtcV8JI4n61i
vesZlUI5WhRsZXZuBLEQDY34bqGU/Hwo6hVD5SrmAAUoukceCHZ5utrW/kgilJ8dZtfmJU5Zy29I
MVsX95kPUbWTzLqEneO/cAtWHsnKtTkNID5YFz8LNbMbZ+WWSA4VO97LsrEWX3iiqko8i2ZcABp5
v6QN5GCCBBVCgNaCyQiKMB3nWmxOwPFlsdDavXHL6LnNQPNdrEFvBhHGn0Vq5KTJ7U+9Eol1q8WP
NuvKHFnwIbwpiDzidt4tGHMMkTOy63zPk3JZJcrRyq6SQ6A5/uXtdYewdgNx3XHtwYXGF56Nu189
z3mgkftOXgOR5wgsksSxf7prxV2VSbP+bJjhx6CHYv29dTMrH8tBhMBh+s4fnq8Ha5PidQm04Y94
PP/4LnsSom5ZY+uhGtYiOxDTtFW5qHeYwGEESRTpF06d4lugeeqx5Rt10YFDaSVkZXJ9A0Apmx9b
74eC/bW84msDVfP1Mj/xVn/GLGGJTVka0uPzIWf2Okq5deRhaOlKTYDyCTezl0cjXPNWhzZEprDS
gi1Xuf3qJGN0sxCmtLZpCYKNdDFER9uY0lgQx9g9AhkelZ6dThdqjUeX17B4p05v6t2xqQowOoJO
8TxifZnxRCi5H99DgcNuAVGMi1RRTPew6oXUYhLu9TRhYX2T9oacE4vYF9JXE8UGoTtJ7jf1J4Il
gcMFOmDRq1rShyyVYV3/swkb9Uap6X/jEd7u1/8m0ftuJkCMzrB73R9uSebNfq8jH3aTy0VWTTHt
+eZR68lnP1CAYnoKE13GcOY1CM472cJw7cir+lAcMYpisrDvWHab1VozzI+A86UsMbjInUoejHT6
hBagQFA2N6m/WV+OFiP46o6IKLpAPS+BFz5U90es+IYvTyHQRo7/9oC1/Q9KX1Iou9eVT24QuIpv
pvf1nJ0I6RHONfnz3HynaPGP7PUfHopHIFbPhNbKSkGDoT2RCwZMboGMmIoRSJPLvjqL76IN9yhC
r+n2eZUeSO53euJpAUZ4A7oUJ1GKRBn2rU23d+EfTS1kmNOVI3OBEQu8sC0sRsELekHkw3KL0Q+2
VelttnhaBkEvS0cmtkbUWIFiJToEkSq8lYPqqLKPb6uR0LfO3rOkJ7hcKdpeN9DIqkTZ+CnvGYEk
xtJnAI3AYhQqcmFwK80VsLxEnnfOB2ZjwEM9kbRgNGOGvTEo/THegONYPUuNHfjZz0F2l5EqHIGW
oeiE4Ub/Qv+014aPSyua+CLtpdkdKLsnIHEcAqhIvAGhyZsr78bMaUQNKpGwvslsGP7rNsxJTtU3
RYZA1PJ23QI4hPjfx1N80Uq/R/L4rb1WzVxDQcNVtUQaaVogv11L/ERMWtL8GjvqHosMa+HCUEVM
iwo6OnNdUSN7/Ws+p9iKWMbh6ZYf/LbZ/rSsMAD8lxSxPzLDm+Hw4jZaFktzejB3cVhWAFUHzJuj
T+QsJxtSOokXCIPBsxnLIpb9Yz85UeBmhIDMKq8+rsftg5Z4TsCo9ZlNkq2Hj086z/XCsDFuMDbb
vM2013y4WvICxzMgQLrc3PTBIb0gsrsZTGsjoGJdjk3za+eK4ieZEpc5pb8FWCTlSNnGbMrerrDx
/Nuynb+R3kww6tJV3DPJuMTCmKsLDTEQdXbcF09Gfm2VFUpVW6RnnmEA2n5fRekxlJ0LOFku1pag
CfB+ucSggh3ZLmt4HhHAB5soyPZCZ8D8rQXFtrtjd+bijf0qsdLaec2x1sfS0mzlIpA8sb1nqJur
QYGF94A+rNG9oKJnDVF6afoR/qFGle0ulwJIBBEKM7G8DxAJYcyyh6tjpxbqvtqhPnMZuoi3lCBl
M8ZM2buSRObh3ufWcfGy1sE9giWA5Ctpp0s2MdLybwO3gKudqiTJ27cdxFRi32c2E4AnHdHDjwso
wtirVvvsIbOOkkk8OqBrX+mKJJVe+tm5+Kw/FbHdYoFPHMvdaZWvodhNeGoC4P7wNxcURRUqPksN
c5GWcy2DHheMwiXVrNjKu5HxreYwpx5gihQJzCJqVt7oFHlANl7nHyCjUuU79PyfQSRO19CDM3Jo
VtEMmkdIi0Fhspe4b0x8ZJFt68ue8elh0OP/U/CTF6iD9ifB75R8V80DoFjsgsHgvCGY0seidtLy
m3IqByvqRGqaNYWfitTsbGZo0Ziiiis/3wfTbhUoV4wO6T8AbC7CkMuxnitJRIAD+eTzjAK7zCdf
Of88hdV3/mGeJLRRwLdjTSn0Q/lW/mFv4xP0ovbNXp0QfK0R2tjodIec5tYe5+XV3owm0GutgrL1
SiqabByztv1V7nN7Z9aPlLI+9hU2BIi1Sc2rW7cjdnESHSdgdEmkDHvIQkpVpR0u8wCd1X+6WvN/
eCX56aXGe629Xq/N6L/+fQF5qZGwyAfKaXu4zqIVrX5Xfw/IEeT32RWZjwPiFQIvOkDa8MMfIjG1
R1a0WzZs3kJCZGKeZY5xq/NVy1IZjtBEdgA+bS/fopoXpOUhoRBs9rdCCwG2Y7NjzM/DyH7xTati
kdvif32fIvC9YCe5uta9EFFFVG4OgbVxBSbM4h//g3KPyzoCYGc10Bsha3Xz4998jpvuAZNCqveT
lL2hy/qIqwe61JfIdMvWIc0EJns+CfBP+Fjqj8tSzLWdk+UHun4JScRd0me/2YgeTsqw1b2g6aE0
zQrFXF53QD3+vRD8UiVdaZulvtYJj3nNbNalB7VfV5T4C9Pg/4zGgjMXfudIZ+KJAk8lR70//o+X
T74yBAqFYpi4a5iUJ9HB7joWDixpAP7QRNBckSfV5TebUIxH7Z3oaPZEZfT/F/YDxDxf3I2MH+01
XVRA8Rfauu5H56w8LcC3EVTdc3NBU6s5D01f7X5x20I9hD7texz7vymQLELW9j79FgNgfMvYDJWr
GUfCTLZ+CMZLIyN3WJKmsNQyTxskfpe4pj6TUN5cQoVtc0ME/QaLGpxKNQD/C5jZjVqY9Z1EInJi
k6aV2s/towCPaekJiaieBPhCpFY/0nGhA7aWBFnNn9KKa7iaWIBLBYvoMoM9gpeZ4fAjvjCYSRlz
2c+upoLVCdgOYD4ThBLCoPgDzsoi7L6dDEsZf4usvI+NO5XEgrhyRSmm947D7ktRBveyXSPNrIJ5
j0VqfhxCumhd/wJHMDJ/gpMW8LnlBfjprMFzB+Zy7+xcAFxWfcoBrzH3FzCHS1eS9tHHTJTn/kvG
eLHRmtbuBG98Mq+IQx64ZqKc245E3PSM9PGcOIC8sTzw0I8Hp8bXGWYnunsv/n4mRZkG/j8iyVeu
IqOYBzG/UcmWotCIayrY+EzZKNjfFnA/gMOctUU0MRbGdUR1Zi6Q4vCJrEp+yYeHS3DCUdrfQpDq
Td+G71XPgZVz5SHPTwa1JDdm8GvjHPLNoBbhz0nLkK2qXTmUWI8w21vn3QUyYwcUBVL5P7MU1Wui
/VOe2td3G1eR1ARJNSqn+hvdGpwfYTKe39gub9qdrKggSl2Lf7jnQwMGAy9pHgP3g2Rlz1Z4XVkP
c5mDzm41s4YtAQHAPZuMNxZU3qOaq2TWgZNlkb5fKIYShLWCzqAKAXuWgyEsWgFKhxqJsRD9lF+m
A9R+2n0h9lblgqGJsjbtDaIeQfhm3Io/yNPJa7x8Ta/uhRkCchyPUqCpTRTTwXTNQh0cbwkGOBII
909Ar3N6kWvCsFgPNRvm20UmFokA/yh851L0F60jcVxEjNuC8PMwAPSO8CK2jomdce5oZ/zYgYCm
OBkbCnUwZgvQiFn0lW910GSMZ7jBxM9Yay38LMxtqWzKVNo4iLpNGUQxVjINE1qP31JJpfbhfpWk
Zqum8OCwmSOk43g6aqZLWhGRYG7xxbyvV6QwS2OvZNLMoKPlxrds56o7iMpJD+TqKFrklaALsoMy
dmrbp0tZWRIFz4Ud1Dou8rrsXYkQHlRDKvOpJszknpTwMYt8l96dzwdh5nnUFYpsudwyRXHJuYFu
gFv/CjJ71I8IXUbvjq+/k85RgEfJ1frGjfXeGVwRdfTKvf9BkW/AoOhjsF130SVnscH4N8eqG5d9
LDFwi2S3/W5QQnMzDnGTbXaLljIiwLfGuoVg2lPp/z3SBdLW/Q3U7O1zhgptP6RCo5YjGZBu+mTn
82XEIVY/WftBV8vPafK3v1Q0knnZXcVhOPs8cmxCpdjyTidndGBdAOTUntXljZpDstElqaY/Oqha
IxeJGBXhl7CllH2mxp6ImUnqz6W38IuvtvPjof99ZUTC+XDJvrjqjEkPzsWuy8my58WXV1UjfX1N
6s1rxbPShf8tajo2FE4tonEIk2juWD1uY4M4DgzM2S4mx18GK4mMQh9M4lgN1zTu6yLbkA6Z+1cj
EcYriVadQxU0ZvButxMPAddlHry/NZpmd7E5aSm2utkTwzJWzeJ3KoI56plAC/qLEkI3osNdDygO
HZwP3lrIA7fTS3BLs6v7/2QjrpuabWTCBgXlAUYXxLFODnlB6ylOYQeleIwo/PMRKQtI5l1GDKnS
lYseu0KM9GF+eZyruJLZ+MukpRmGiHqFTM4FylNWwxuweDUB0VzOxEoTsPiDkkhoKMKNuNo7okem
zyU5FAoJImBiR2u0zji4cGxbmc9cWCbhO55AQIaWcszNUUomBMjmVqjAedSQ3sOebJfqPEpHtizl
kGwbuHjSxJDeicMzz+RjuBCAA4qO8NyorhlZxvCpgg/USu4/UDOcw4cckyY/XJzAGN+wvCEoFAxR
GbaaJrjFxl8Y9tUNNKtjbpwW3jpeHdC5EdAM5XQIIUN+rk91m91522TALY3P3Z6w4yKZ0izrQIE3
/8dSFMNSjHljfS9CWCJn1XE22OCBfbNKOz3E/IKbwt/EF7Kc3u/rgiGfCfhPVDxG1j7dgMiHwIX2
HKa+/PEdDcZ9kKxCWgdhE0K738H/bSwfiSjPsm04mLpJnbd6Wl3ozl93Anmuqx81yd5s0wZEO3DC
l4m4pPssKZ8MIBWTnYAE0vC7kn5z/9UNEzTLEu4BkVpp+OlgKM2C0sxXTREu9voHzGC0ziiGZNZl
HkedQtHdyQk8DkJf5dHE57e6C3YGcV2NokfDbzcqSSaUMXZq1bL2MHuuOeXssbAMlJlJDFyeyPvd
WGj0P5Z0BfVPBskEWg3P1jq6mN8Brlss7PtwNWas7rFSgPJdowtxa0Nw2ETyf4AL/W0IUpxhMjN1
hE6j55a+cDFRxv+MkOeYY+rGNBaKqtucGOD5b41fbKVRCxo8qLupBcJOSy/MJzrcmX6E/sXyQhwp
DFeKTKRSnBGpjvIapbAAKTlmFhSuWbXk1VZZW12zR28rsu7K+WlZYHggxhY3x359gYBILpiDQ0b6
hK+UYHxCJO7/9+EHLs8c9v1G1HvF+PziyOEARSc2mUeTi6j626733qO9D8XzIbMOZrmzrQESNaCD
0+5aywv2gMALbsvBX9OQLYlOPfh/oS3mUzBqwEmc2Kgvj4byghgviy7yqnFayG9igv+nI0Rsddvz
6C0pj7OxUBMqu0MIupfjEjkbhYJiBK+k1FP2/fZ+SGghxRqa5CrqM4jqQVEZw8SJx9rgPwOY92Eo
nF1cbHW3qX4qd0fMnJl4Tq4QUgNHJ8KXs99LGhqHgeGK74nkw2pFzv860H5abChmrp2UCrCpBsX8
3zqtgj+uF5H2zneI4tw0Ghm2ZvsALDOz0F+F3nDSpNnvGweupEM1PJVhyjWqpB+M9amcX0wMdb7+
wYUpd6zklemsCtp0EUnIEbJDy6rpol2JXPHBcSnX0Rc6EPY83cDVz8JhGmCFX1WvL1iaDrpFy45X
lA61Na5uSqZces3giFl8vgcY9dGkn+zfIZ2ADXxy0S59YCOpNWiDstvSGWinQ6ZBcLwsysaBuouo
AbCMz/LpTPij8NNbbm6AixE9Kn8+qWXxHdxFS190DKy4OzTLqT2Hes3u5+e909RhxA2AIVr0THxM
URs/wf8CRocG6Zj/JZba1GQtYhIM48kuiDNAmO8d6NHm+ZvWgqnzZ/boizG2KFqBXvAkQpKRrtOD
Q0JkEwFtlwWV+pP0hbsFxzaQX3uU37rC0GKVbtsr7I5d3aaekDLwJ1GApgdg4AZPP9rNdbqc64CN
4H9t7FhBxEuIeeFikKg3v8ZWrwCQn5T7srIQ6tu7AiClbMxckQVn5/r5CLLmuuvMTkMqT+6UMz5M
XFe33nRTtev0S+bIdD3KPs/Jc2T0NkSxhnjcBbRUC35VXligJcF6Fqhw3V5g5nLn6wWeiR8xZxn2
/Jk4q8ZkYxlkNRkonjE194PIWDl5H/5VKBUz42s1jUJtUiQyOdjrbrj/n4kw/3vyz+wi3uvDxLBU
50t3h5SVHPWc3stF2mMB06wR7LDtHG5eqhGzlJd1YPDPbrQRXT8qE7YaCn7ITD0vwTTWLO7ltfqZ
NfanDY0jBAO4YEoaei5jCP74X7H91NO1RKUWX8KeL9azriy8ITfSzieLv0DEnlIs//Twi5RV+j7Q
nrQgbgrvIvYATxqoiNrhQdvdN1Nz/oQ9FZ8pdC6k2yHh8vfd1hnopnQ3LF3k0TLtES1AA086XgaH
LR6dZ+6hrbTMpIn/VqI9dwv74deGqxH1LK6AENwhiW7e06fElGhpObEBsDF16FX89zEdXBoNy/j/
MuWZ99ljIc8WAvW5E8mBBBMEj779TzFhmL6Er9EXXSwbuxrEzEORsf/BOGNqmljbqD32MyZvIWq1
Cpp96Yh8YnhVQ4oZO9VdBd59LYUEI8q+O1YKIBpNLzaVqMyn2X4z3iNMowTlos5rLt18ke2eUJty
H9SN116K0VV+Ebi+kTDhGoAGPGxXkG507WmDV/Wn4NgAReDqxhxIO7qetDa3tQibZKZ7NeHhyBv/
0sGgBIPcauXgkVMM/KCUVA0AOEudkpESVEx9fzOAmqjJJKhhhWaqJBwbf4xG8MLQh1EMvTDzdBWE
CtkfshmCj5/uPko0LjlExEXw0Dtzmfa0rB3ZMQjQUnyhtUr566XjaPoBI4BYwKA18h/qiARquev0
/YmRqN7/hsJ1PamuDQfPeZZFBaRN6kLixh/mLiV+++CjBZFjY8h0592nS3Gk9aNidPV+UA9Hdd8z
lx4r/SquEEw1mWXk4IQGEPNAvL9RZioWY8y1TuenrICH3XoNz0de0RqOhp3wrFYghdwC99TUCvpp
TV8IACdGEZIe+cwFG3jRWP3l11vNryG1sAIl/8emgIpAec2rRTReujyq9vsl9TOOt7WK/8VjlG3r
4m89WWRHviXJnipSrOPIS+EBcxXNoDl4yzZQw9wKDphoJq/fj/MM9B2YVKaOfpIy40XivnsneQI7
uqvqCgv5bb/Gihw8fIZmy81WIPJMtmtLPVIe878QmpFXzcInPQWSKszhYNYonCsAkfy+IAyww0ro
MMfV+q3HEDizp1OvUqr1c7rTbllYbnRcuE3jBucZtg==
`protect end_protected
