`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VqeGAnaZK8woxnZL8Z2YZ6TG0lz5tP8zv9PY4dGZUVJgsH95n36Gsv+/I6PuYKbJcv6A/L35Une+
RmXERhDFzA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NeCSFszNIYwBF/yleqUDVFH+VMa59fg4Uvk2VRQ0w0qB6YLCNe7K+lD/1Fm34IxH8FzR5Uwx6Xeg
JBfcsLLeTXWLYl6CP3ZNB1TvVWLlskEkDPp+TB3//bCxyP9lbtUOH8U6/hjGjCX/ur2SeMvknUT/
S5ty0nEUGCSGSI+ChLE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u+y/6/zWyAkR1Tce0J+SuawEEcHYmsjLICc9xVk5CLf2o28EilMIMu+JPPP0Ga4KG446yoYQ0+lI
bDoaLU2z6EN/UHXQX9wCxIp/xs/NQhK3/ztmRBYPquWZ9eqdkUxPrfCHg3ctfsE9qn3mfYAjHuy6
dBnLM6FMXmPe6DnHd4h37A1EyoflfPJ63tWjf6jrqElh1vVDRS8Skmd5lP3Im9jQLSJdnr/QCHcb
iFbMdZ+PGMVsLOSKIcvZxpDlGEt5tZflDvrDqymAU1HwNNhpSvOU9YmdSeM/HTC4VPqx4O6qk91A
tGO9xBKkrIZVFX7WN4aXT8wOxTTRBliE+tythA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jsHN06oPSkQ2UVaUKWCMLRviRr41a+6fMRvTt/aJ46ChiARgL52ph1kU9/k642INXcThJJJxEH3C
R9v/nahHoPB0Ehea1q8oS3ob71JpqqCE0K990vpAcJxdbjK8gp+DtYH0CazBxSshGbbCvzBCtzMR
L4I4KAtN0CGzLD1kc3KD3QI1oNHrH/mSox1DGFShJQfm22IsVcXOYvdon6H3UjN2ee+x3KAO8+M8
4Apvn1EhvKXMS96B3DgFCDQWpXqueXXv3TmBgrcIiBRPnaq9ivUnCRG5/TgBwvFCo4b+i81jYP25
ZyJTJPWUym1EonldP/ueH74gKpkn2nNazYvovw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g5pddxFhXDVpZ0YhYmluRwZvpJO2aSNPGGO05oaGXehLD6q9rx5og+9bonultNarszZggAghmky+
8Whj606ytkiFus4hNIt12fmHCDub1hiFMO1uxCWi7j4Th5mic1chtMyzNeIaqTkTNK4kAcJsoMRv
LdXKmgIJYxWAGaJ1Qk4uh+cza2e15TZOTGm3KCEWo4bLFPvg0d4btXONP4sSrbQh9XiTkCibszYH
FtPAqY19HtFb5WNdE4TA0mcDvzWF0asUGV9WMQd4ELmgIrmrHk+h5cDk9JuHMEoyQiFW0xew+vey
gC4RmWsZQ9iQ++Kp5XIIjN02UKh4TPsSStXRUQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n3RgHkmaSwLLgk1QlK8GZqcsYi3QWmu3ZppU6kvBEsUcVEYkeXnWGRtprr+fofDe0vOL55U1aj+u
1ZNHJLa3iJd+jZEJyazP6zgUu0nAM3MHXI8Qol72Gy8HnYlnf4I95pFTZCUuLTMSBN6OgH8x5yGS
nTAu3azVF3NMRKdyw90=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WTY0CG4JfiD15nWbEwTte/9NQ3of/VE3j43Um1mNm9dbaX/EbcRKqAmmA1H2UPmK506531Ow0hPn
ykcobkelSchL2udh2sOMlRVkRuOpc/t2JbFw0EHmml8yfCNbwss+jlEEgGwN708HfMb1v30nl04b
5qoRHSXuwUkYs5++Zbu0z15dmr6RBddmUQRYtRnWavE9PWE4yGBSXsBPpYc/7fXRmStqMmgHQU4e
2bnFns9AGisdsPamJtQdevj9IPqddUvzsSavEpZbmuoRlhZ/1ZLmmGk+QH6Y0n27y9owVumISrTy
lDhD3YRNqxNfpgOn57pymJsAjCfr98XqkcktQQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99632)
`protect data_block
R4ZtrvilN7XiT/VmXznPcp/NO6GylDmdwuTtpgWfcA8kRJT4CWmOQqckBh41wC4zHkj3f9h7mVls
NJ5H00+NkEebh/DWd8ddRUAVUfcGQ86BcITY3+dwCorFu1/vncf0DLazSsiZ9/uBpMFqralVOIyb
ge6V7/E0N1VObtazFqMHnzNxRGRqiSv8oMIn0XL1MIKCIEnbzbI/fIJVjGdD/w0dc6TqKVybjOT/
Ld0ey0kD7jMGAbjRUvpTiQ6q78INncprBEDpe3JFOrGHYiLG/4Q3r7w1bDMuudXqK+XFbVEM/SzW
seT5z88D3ZQZE+rRFxRmwgpDfPNYlsCdg740Ofr5sMIaB64/jOWd5Axfji/2Dm4lroK+EccLO9Wt
Z6nP7i2iDXI6LroCe+TeOtomjyYdVWlU2RNVx/IRmdvlltULLdrfdqyYv3LtRCubC7wyV7532QS3
CDOv6rJ+cB2HFppztqYkCJ+tMohA4Gw3/onUAhzWAYZ645vPDEPe0zgFn1KWyYYLE+yDAgm6mFIr
ids87zfuQnwkVpzHzxGfkvxPuTij/2oYPChg4UR5qiKMVuDPqKc9u0yvlGO9P+zHZQEqgiLrm2A4
NFPDjiqpGBv2dlchzjXtPxWos3S7S/6JbKXPht/wHRgjUn3qWzVKAWz+eGcogaZdB9G1jbBXmZOF
rPvnUUBuaWkiyAW11TBZcwR6ug0Ganz3miD5reKmJvZYXdL+KBmUo6qRw7Eo3VnLUMjPBbjTKOHl
pTBJLX0cZP8S70eZJdPRagIRr982Q+O7AdNEPZcBXXkPS8duNjzY0VGBfj3891r+ECgTZa1gDMXe
vJDoiXWVklasy8vk+KpEbiugevRd/EIPKssV/KRD86X7ovCZ1aZ9JouT2Ehy5/M9JEcFZ7dlprFp
yBD/4e0JhqsQCe6BcHBlrdA1WmOUuWGHV2ubvsu+d+fErm83ORWYE1buYbtJoEAg3oSusf5Yuuik
5/2zDHmCojFUkSM+fhoHfduSZ49y4tOColfvKar+B56a4PJvCs/4wGdAAID35PiLOlVBJ0LI7E/B
1OcT7vCJoDv+lxg7IZ8v++GhTWiMK8omGvlMGl+AkgCkU84Hlroa3Fn7/NLck2zcZnK57TNlegdH
fz2ayYq+eEIuGJXWEx6S+dpDK3W4CZpqoCwX5+l2PGpHGKhOqMII86uz6lO+fF5oIGQm7yg71xT0
BHOvR8ujL0zLBm54YRoM2gO32zVqJ+QBgpKyDC8xOEcHgT6BI/mAYWP6Ml18pkmITjd/AiYM6Lb3
8vZHyCvXgM+bzPF/brhTsTvRVqQxMOu+mvhnASGjiLG6z6EWjNoJ6uUq+wgCdIhSbsHQyIOElFYJ
bCz/U0ZjRby1cuMEOoKhG4ZPfdPu3gt02D5SzU8QUqpEyKQ7YeNLz+48S2+tnOvB116XAL++5tLy
Bmfi+9qVILd29WRW5YH3Lyx/ziWvS3DFcSJaJr6tJfdNt5aodhx0h617yfLR0Q0Blvo1qnSKm7pL
WPnQTjZYdQe9FVxrhiBBBlxNSj66FvIfyCC1p4Kc4qo+faBoKNVkkpqvIu0ukyAxnrFtsqkdW57S
qN53YTP0hk2YKzk0QBlaKsMPROy4kZjaHJleReWHROWEObRYRqFMp011Dm81xPBXMtsEZ4wrRwNd
T24jCg77L5laPjJXuEpVCFwKYOTFXlc3MdgzbSWHFx0HhnzVMGAvLsa6vUR7Xnnpu2bWYOiftgBT
HYg2ir6wA1NrSxeaqOdcMlQ+tfwB1WvERRL0UuDIuyT1oD3BoEVsibXBznuWac1KNWFB4sWxUtSU
z4/njNMqBvzxwSwdGOGanTI746jgueoj0bDsPIdOccaPNOGQ3GgSgqyyzfR/ASZL+0ijnEYaWnmv
vfXiJZGokFea7Yl83iZaPW8vzOjRKPufCmX6YBX5vPmvcTBGfJS9EI9HeW53/wm1l3RkgPSSut7o
/54tQLbDYz91WWfHhAUllVqOBlVItvzp6mKav+ZnoxlYR7K0ggRLlfBMGaj2PJWWtv1dTtiMWtT0
Y02UZoBA6MpMZ33oqfjzMDFDC1x0I0SZ3ztiv9HhUh6+FaNHgilrN2xGsWCK9vvxJWMUQwl4+rrP
IF0P2g7n2klN97qbiZjZ6xKBVsP3WjZEXLNFJXS1HnZcnXE0IFlStj6bYojCaPUgSSnjTWyzQLUr
X5W2pTa5qkCe4mCrMWRkvRADUzPbn4Rzkx0MY8GH8yff5mG3qp0wFYaRZai547sc6S6w9RB18A7G
2XvpHQZ8b89kiDL6cY02Gl5wfnMWbHKjZTg69sgy+iXp8AriSk1OGlDeDp91fDuZj+zqFna8eiOl
lpik/xT3MUd7zO6jc9LOlhHwT1YejyrWm3eg4HlQ+CsNpFr7J/v9qenq2GiVx9wSLYYSRl/5N5EV
ihcWD+dEqXO3GXXDwiKXeQ7zCNvtC+hCMLoDX80e9CBKfMweNBmvlkgwr1MCrSx0yZ/KtL2FFV4c
ICXdVUC/CdubIvGlhTh2p5kIurwMqMl0qN5iA2L1uHHQ1REFzlL8HkxMKU0N/E/lMEQH0+Fn458Q
xUw58FSQtNeoSvF2ZkpJ8brYQVSWQpaf5nUIqYimY71h2RYIMP3ziUwimhVCMT8Zs2lvAHB7bLck
SwCFRWR4+4QYStBLqi1nRPLGsHjD4uf9eFJJJoDW5rPJ7XbrYUvecrJswtEB1+NNL0QGa8IdYnbr
MCIWHIZBXJiayLgoX+h6VfDzkvw4H6ixZW1XiXxhkXGpgoz4RArv9uE/a5XPz9UbHMRQYODlNyO3
jFXFf9h8YMBVQHslErwmfD4df7+DsFtWDMh1xMK7Ixe1tAyD4v+AIYIiQ7gWGF9Iz/Nf3BXjrRz3
ZHKWYrpJk1SOGTAQW4YGuc86bd3MYxaqwAKa3oRz9ywHLR4jPgw7grSoZkCIS/dJ1galT9cpLGNr
EFq9fMxc/sLnSMZZ0RLdtlBuTF7b1avZHdlQt85IszOsuO4agjUaqaVX8ZOSAyXqPY2WeoBNjj5R
AqErNbNYQX66S0QomRcZBaBVp0jAhOb6rGdIfzNixmELra0d5TClMmG+bi6uBW8WfhLIJ/A3pyXA
mHipXdaQJDcD7kq6QEeXUgsTgO4t4LVRv/qt6LUDHIHmc6yRw2O31DWlpFM3lN6yoRppqr2zx1YB
kTnAX7MQCYUNzqsmctZV2Js5f5A34u27aDXda4BORYiW/XM0O26UlF7TtISibaOCUFKgNxtEoe51
pSeD48JmSd7Dw1WxLUJV9ENqDAmfEdi2H4nZSWViLq0zxe4PUnf11e1/5M1VM1f0FcExmiqz/1Ew
njplDvf8Pfb3kIPqXTXcpI2EjhRK5tvODDUhNL09kitZahrcgFXfgVciQfji5Y+iH6fJDr6mOr2d
dEgVamumHL7gEwNxMtjwgkjECls9+E9mYLeRhD6tshIzZDyHpB29sgpemka2ZVCRgNqqsmaVu8Tp
nUYPoQGBhrMz7lagfthUBMtEC2ghAdHwDY9WXGfNyr7BHfzce09o8/Aecxuqsl5qjNDE6BW2LkUR
eVZCfnIUgsEq0OI5gzCJhcK4SLWKdei9rYqvoE6PdVyJXq8ht/sk17fyy+yew98ZRx6pWBt0IAc8
q+xaHa8KF3FLZaH7eIbfPmjX8EM4RaLxerFzQD+kbYabZYAhIkTS4rhGlPjcd+PoVnZ96lx9HhG0
n1pxTeViogQuSyurt+ClQCjMdY0cW7lj1ZTXMi2Lzo5tfIrBVFZ3HTwfPVJnQ0/DoYwY1KxLYsgD
UxU7Y/EKtMH42AOatn/W2ckCNHlYUUrJQJtl9ZbMRF4x8EH7on18KDISASwdpY6hwikOa6VnBtAB
hqW1F7r7DIjQAMuSJM2wxZ9kjAfGJDF2xurn9jKsmSC+rjuk6SN/WCpqpI70VkSV4OjMz6xxug/j
N3jwvOqnERjM8y5tmGp1okIaOR2ZWSZq5Jav9iI/CMOxWHG57AuomQIoVCoCdfopS1e5Upz05rL2
SqduN4plV8yM4bgDwgm9BNS2VxRatPhWlbMo037iCwMi4P5slVZNjhh07wfc6N3U7BeSb3OjzZHU
ji7eJHiMWYlq7+SOXh6tGZKbAyD1fhcgsk5nXb4Siiv6xQZTopt2ejitW2tzD38KDKMD4T0Tk5Cf
ur+okMEbQBbqUZWdg6IMwbFNiG30eqbIUGc1pfsmNfnR9r/WDL73DOr3miOV+wV/yjwOMWOp4GFC
fHJRB/d5Qw4tWrSseupqY5JWWSByAnHVJSqVJgw8E1wgiXcMAnKW9N/4pDUPyI4ELo1+km0zANxW
T6xQF+v3rM0gAejUuxITkvoHZYlfEbVILGNqJtjzy9iKih3CfsEBYxjK20vikBO8dJyuvtJXRb6u
PsSJx0EcTVEoZgPSYjFW/w0vN8UXOB1nApGqnZ5GKHEUhtcZ10GWlH6YT2Mon+lHiSubO4hNyjJf
2TwrQkXbFKn8KYWIbX2+C/f1RYI7jyyLYuwcRglSg9nYr8gsh4wOtTqkqmYGnaezyzHha+1wjct4
08FnJ8H7EKoWX164TZCxDd2rkq3nG66xf/NhlK8AENSn2zYpdEjvRcSbTv/HmOma77BRX61930HY
FzPeIwZZlZp9cv8eI8r7FOz4/ZiL5Um5OXgW9XbD9SePIiN1SUH5Wmk95IU3/1RNN4LlioIyz+qB
x0epewuLNTGkaLES8a7iLAkK1sGhRGc+4/6k5X95Ft2G067M/unqKVUu/SDnUsCqQJIRNlTvniFv
ppjL7jBimOqTQeZI/NA5qQ2NnUkE8G4oyQ6EguvAnpsnh0KfsS9Ic1HfoV1aQhHDTGnQ9UJdZcbo
oB8rXQoRcc01E/W4EkJ12S+zU44hNoOFwa0ZxSJP0tSp3gKZZoc6auN25z8vULcLVVHId5w0T1EX
fMsOqBWWbrLf9Etvzx5i1oHtwFyqE+8t7koJXSHoN4Euzd26y9Z6jWkOzsrG913FiViBE2qYdSGv
5J9nZfLQPu7khq3IxbKFZxQrt/db414gYi8iBM+4p8fqXfbvoTX37ZmgSBmFXElMAOoEj2n8k7N1
rYkb5kDq6BQIdgk4zNNhKTA2eIwsp6yEBn+f/YUYuvWEyHd+IB0RD5Gsxye5SOV1Ug77olCG9Q7W
5CBuIdVvGmHoGpwevaAF8emBbLGlZWLKKq9UsUUHWWcJ6Lvmpz8ufRMvj9C1hy9Ix1UmK2cy7VQ5
5dsxjcFNu6KRCMJduF1BIcbWL23XPQQTV4G+Hnce4XD0+DrVZUZbYgfNtm3MYjQYecjyyPTZjGrJ
fDXQfR5DbmIsls+UVh+07RjH1153v2uqWPsjxhGNcb8VxBSA3m014agNwyaDpMDAolH+lJNaIgoy
vgXA9cj33wBZJPVb2B9ffWu8rf5x8aPVo8VgWEnY80eu+JGDb3vUYXYvBpHTAftnKMxXhORzJDJY
PrqdPSN0Ozs1aFtI5aFMgostg4EVps1yhfQoUtwfpMprwQloPyTHs14DWNNLpHnIm1dbyCG/pdD7
MtWqKx89jAyc6puaq4/+eBJUgvmBHvTxi2g5t5NCnXHxYFsZHNYB8cPI02ngrcVtcIDgp6xkvhZv
I4mNk1cM6kaPEF7oIjuWKI0wsqc8LBIbmLu+IF/hWBSOX5ZhsG9KNldmfd+Xkk4G/aNDGz3mzoi+
2/bDfEcEJSrAeDOvzKEiYxpXrvhpj+4ywny061x69zv2EdKpR0q3Yg3dNOXQDSMdzkgyT8l2nBF/
z91vxUrN09SQlCUSwmT7nwcxRg63gXHUivK9MgSTAPWGKMurkx1UCknTzCf2NPOPhqKIjz8N/tLJ
eiyDRMIc8oSbjZ2cEajsbHy51hETx7AO4L9G1Q+nzXvixFY3sLUbLmv8kZd4vTrry2a9kTDaKuZf
YX50Yxcd1ez7VoYS4WrOrEaSHziCEF7PbDJg4dmEC0bqrdNFt5+suScNMCjKMTEHfrXm0ykv1rnO
dP8YilCUqYZC5CenIQun05+gr3xUfj6zT/tZOgoSzp1loBc6wn436zFQCi5FMS6lAajCtNqAcYfB
qWslJ0Tlh1dbeVQr356iugUeY5GbCFKOiFp9Nt84+dYXPYJYkrTy/y/gYp5saoq0rxl6kkHp5qzF
xynXBzbBv+mluh0cMNVjN9/24tGASabbF7G+qpzcl7u/mNxkoIXyTK8CX1+aYipD+KzNOMmaoQZX
0UmITFrWzmFgX2FWBL+hy1AK4kEQ79cgAGnXc1oO9h7gC/74JXK1TM6ecHfQP6S3uX3Y7d3RCCJm
oRTEzN26h+vS48fbYv0S5ZI79hyhOmgoWkOV+37jlJTPrfUy69avmhBS4gqjoLAGuBaP+vUqRAnk
sReQFBkujYGZ2NkrO1UIVK5brKNIUhBmt2YmLY3/V1DOt5nKFLtkiuVMQgIdg3n/GooYT7B8ZibE
Ik2ZZ8cGAdK5JBiN8aSus7Rnk35FJ4EJSYtpeMhOl7GBKD8/+EB1ljcHcQ3THnHRXpGFyM8RQsx7
iCjG7SAerXK/OntxAJFrDp5Llr+MrTG9eiM/B8ZfGXH/9XwKZJXJLq9hMe56HsQqjDEc4AOlVLfE
TmJNo/wYqddkXopatu5H3UGovTq1au03RjK1SDU3TJnhMuHKu4cvC9n1H8rRtWLM/OU/DpiVMfD/
qHWs1JD7VTyiwry+hBFpIWEjpAdh52L718wz0AlI61dHE7fdK/FaUdJgyvlvB5ttpd0vwUsfxpbp
r5oTvKGpUZWZsOER8aFbA0M+JFlcZ2Xy7QHEf9+gLc6GOPEircfksFaqyj8ff18jjg/cLi7A59ID
r4k+1Qi9jmPvcdkBZIzmJljCUHdRNW6Ceccb50s3ESs7xI1FlS77lw1V5+ABikZJtHEWeR4qbpEz
fsn6Lc/g9zoXuIFT1JTQX2DeRe3itCSThNTOeICrXHdtl5sL8w11Xq5gfrFSAvihT25pNPolaQ7k
DXI0ZuowLLCDzfi0vpGHKlRKkLs/xOV65CVtfEO7h14hhbIvtq3G8POEvPboWOAaRbTQiLnDEwVC
9AjhKUJmBAiIlEy/rm9DfTtqCIbRCrWbQxTsaTX/6BoDbmK0OtY8ZWSUYJd5a64g4Nl7XPRTRCTG
MIGuPRPemuI6I5qwWpn7AuXlyeFGHYFE4qpXpy+PG7wDFIOr3fDYrvAWGUiHwkHEUkp45KQFufh1
YagnODAiq3cGT+5G8gCEomMhoeirG4/Fnzb/Ce0hwM2RntQdaS/uGnniTkt5RPScykxHDqtHMvvp
0w2mZICAa9qGrua2LEsJpjd0Ga/QC4ug93XT15H5/08VJGK61vu79IYvy4VxLGn8ODwkuoFQtv6P
RjE83P4Gx/Z3q3dYlivFqr9sgQum/wxC7RRX67w3J6J+LPkA5L9JQpqXmBvLqe7qp9DeZpn+xlou
t9tvB7Dr4sG3wB2C3V7NH/8fbJo1mPVBCVIYaxYRnpSvzlnEkowiUBFp7OLGHgrXLKcOq9mmsGch
FuCgVB5U4sJHH154v6zviNuR8k6ZMuBMNset21AXUKXhG6qFv5ScuZt6X6sA0lQI2TWaN27EHbCF
HOykrjkf0F51I/z5JDMZ88JJYnbNaXiu83j/98gjNcty+F2nB4hzwitIzuiJlnZG8jC8ArOHyogU
PeYMyd7qWM7Yp4zO8iJpk0qeKHwnSA0dom5uxAZn6/C+atIfQMrjRKoVZOt7Ao+VqNN3bDaEy80r
Lwhx+JWtoTmDRv453Qs2T98Vu1bnl6ptaz8gTOrhKiTBxPTDY3BzqJCZIdXNKZunKYoyd/sRMgH2
ayH7CrUXztnRhkef1DH/SQk4kCQkUIiJgyVD3wLJWrxPUTv4QeBO32dw9zTneh4RkQPnkhFgMCmp
OfK0Byf7NCVfDH4f5zSL55v7iEBjElVUoJhEj7pViaxpTP+6cJt/LBW6+3WBN958wBWfx8FDCUNd
bmdvfdiTIdrE7WQHXA91TIT5pEPakzu25IOm5emOowVsAVhswueCzdOiQ8b+KplEb1gqyZ/9dHc/
ehMRCIMS7yDRupe7UbZ6CFwsC5PA/8D4Bt521HJ5sbkYMnV1xuyzLlNoTllcqidELVwFlu23+Hf8
zbbANPEDvq221bZ3ph3URqn28XnzpvmjBYzdS4fa9+ycmKybLwgSwKik7nu+IgLnLS6uaTOZl3uR
rPuFeZioHmfnvYpiIpAwedaMmTtbpMnvSg6o8HapWpcdHGeS5jxG0DG4gvDUZZop7lspWJ1J/xn9
tgB/+1EGKzMhgpnbFPRuQX4y54QGWS5lqm/bA5XDUDRR2nFlW0c1+xjctRFDnXs30gYCsAjyrnb9
Y3ANkS6BmLIzPc5vBaBU/qDN3RotRFMmM+ZdisXzp6p3Qh6oZZHNDnOsfLss/Jyabr6b1tHrTf+p
Q+Xytc8dmbOjEba/Qf2U9vlVW/uxSJ+sEnZyLkLoETKe8swMdvlL3uo9uzPCRkzTbqh61k1KISIQ
fnQhDcuMcbptEBfJ7MzaxTqvm3CAYH2Gq9V5A0c2y8HP6n9rMIptv2k4KVdD9j43s9nrkXVcy81W
st5KZqiDPHvFcaa8v/6HO6Xv9RIVnp55Ax2iN0yEjIWvSFoDhR+5cP0Y5LXgBqsrXnWGDYgM8WHK
0ujFF4xEhzL3tGz57JHFMXuttEFXtt9WgqFOrarvlcON7xEzWw/MYAN4ICSCi8/9PZKEfTEDuxrF
eosjRtkeS0kOdBB9y8MMSb2wr2wtyzom3B7hFnJpq1L+tAIH7rAI6a3jMdFYC/9A8IWycHRLIyq3
HmR1aJTD3JT2oytM7GT41wvSroK1ZLTxonybBfhv6MtOesBb26aIFK8OFYLVjvLAzLamiKDdZgF1
7yJcz+Umvp4CYvEfCNvlOYucWu2dtf0uZ/o2/iSqVhf9dcrMDy7IuQvMV+/IJ6ZAJICFMJ3oM7ZM
QXP1iU+yU43xhtpzEHVE+T1dKQJhf1nQBo/KKeWMccBjQoczusCO5nQ8YxodsZFdBKaKRQ7wi35Y
c5G9Jq3ZfAvvpLcj42FiF95LmEudrIlnZcyanCQjGPFvZTCETIDGlnCIzTV095o9S7Dq5tD6Oyp0
edqdnREWoQeUfau7dxkjd5CPx8FS2rxUnhGjaf1lbCL4PYph5dqH3y1M8Sxn6RqljeFf+1Dntj+O
opKss8KFya4wo1tvsxuHDPwryJSPgJgxIDV37DPDJJXtTCH31BV9AHsqngQyGww14WtYPV1CN2wL
Wh1tJWsPz8EibwFUz2bRdzFkR+dML++L4M78ON32nVDXPE/Nu2k2DJZzhxqimbAtQ1u7D1UD9Oeq
+nlSpGQ5X2owCWXHc86TKROkhlCDIi9nk2uaiBvSZL+MpztWoalQvyOYsdzCxc7MvCkXLDejmVxv
3Mn9m511H/ap325iiZ5ZGHXkX2dZHAZ0bCIUFxcJo0pWC7UyqR3eANlKx+qNOl+sCfSZrp6GG/dL
bmt4Ks48e2QNZ+4tpGalmAqHelBGfhC0RqzNWqPApPEEjJH0hJmv9tKYVtWRwVopA+A8JCV8ikE5
C/8IcLw8ugiDw/fY+P6YpMFu7J9n+a1jjwrzyo96shBb/fq1xeXRsVKUN6Y7YyBmwSlI3v9WqDzE
xF7udUx7x/xcNxl+EBsosNVm9+tAPybrPYsb+nAFpJzc1+tyY5z0VI/jYse56JLGnNrOTXK7i2fX
oj68irvMOoDpololqipKdQDergKTi/iShcR3WYziU2dKLkN4fCE9Ku3mXZPNz0Mzzd8j3k4tK3RO
iCe9ahLPqgJiuvFbRQipOZ8B67fG8w4W7uODBZPfjI39nXlnK0ZeaMEJzg98+UU/54uX1pI2Ysya
OL+xt6y7j965Fng/y1zIxSHe+0WwPjQ95HvFxzFML6wom4unaeAT2RixBeZycrJhTMT9ow9d+z39
ZlDG3dZJn6qp5EEzQSr35TlafbuZLvzeYUnBw8IFKdh2gY4l8UiONSPDhLQB2QtMLv03gA60M9wf
IxfoCf0ui4rkJU4a86wO0SQDpAf4RTIHCg7tqATMXKljk3LEFfcnDabekZlnaziwQpiZ3cWCORp/
1QEiG70MbG2cZTi6whR92g3ZDllptfXAv/5gOu58lun20ZJyw+0h/9heZrMd5NnsGlMQfftUl+zQ
gl4EWVm37TArxB+rZsYMOnuqle53Y34vsOFErfW4+R3mx9ugVymfACnKsrb5J7E4FvLgZAeEI8Mf
veYCzeuPWeI3PqAp1pqw5EDXMGMFWtuu20phbmXEfnLsk/tTzh1PeiUHhJhQcu6+9VCeAgGmM5vM
KeHiPoKy0xvm/jAImwwixnDj8aL3dhByZjD6au6JeChZgR9v9JG/osOdbwhq1hOFTjhX3Y4M0lX+
kgwZCQe3RfD/l6DM6u74A461kJ1fOueLxYpfsJu240HeEzC6LXtz/jiqzzvBt2rgPGZpw+mPNfBY
DDCQ6jwpfCN5b2X7jCE/ZJjxHUuv4ymfI7v21x5AA1zhxdbArXkSUXwed9w50ZKCYTkmMGLOON23
rxjHagJHGjSys2HXZmEOJ2afenAD98xB/5/xRZ1G2O/ueHlGBUR0vQNxgFRlDY0Mggm7isewIhHx
sqjkYxstRWIOz0Q3smCsvR1q33BSwUORuKtwDrdPZVTbULS2ARAppMPLqKX3H9G4MDy6k4iLs0qE
iPVNz+5AJFpajtudr4aMwrp5Dcd81xpO/DcoTU+xEADxFPCZq3NWS2rFiUNIXgw/LU5GPFdib9l0
b65uDYaNRVDYvmNbNJA6d8F7NDxItXTnqf94+UksncqUa1balM3yGgMHI5DNpfsTz8KZ6qGYnbxr
l2YKaSuYxvAjxih1Nfd/2plR3iqaHhrlCINZIHupKD7LhMTG+JVFCiJc7gKfR6ddKQd6YWmbjdIc
uBEFtUef6gVIIl5VBuhxAc2bulO0oftqpHe2MSt83QCOfc/V7bcemmHkbgBsfUnOIWkcW0OINTzo
zCYXxivKs9TvRb50nB/BvtNHxac1cw0/wOxo4oE5GY4fdJe2cgCfFseum/h8n3jHKwM4HE4Cepyl
i4459uLpZwyXUjXfwmD/iiovYDgomsK6YdqqnFZn6nYCvSlZcXoOVOLU88JI2y4X74t4J9KknMgK
mpV60fmzIqxR9naboC19SZveMY+ztA3MYNFM6AFDF6VMgW9A+hae004qDyl4NjZdj/ax8zFHHiuF
hnk+N0MfUBlhOaBrcJp548zoapz+wc3q9Yz/yQlayK0ef6bExnv1GovmPDPTGFFqf0V7waDhfTMq
ugLrJl2ULTnMv0ngjJyE+KUrc/B5s4/bhzwuJagaaiyIZI9RHzX01W+yv9GADor17pa3t+eoF/Fr
1OicFxJo1sRrMZVqo6CNsgWa2/jrFlcePaa5dpO/Nhu3ZW/yQdHf5TvX3lIJXdgwwz1w0mdxZCY/
lbYc/kH8XAEIulz2HejquvSrz8NV8aD0AP/AxRh/ZiKQ3H6Tnyef8jpMWK03RA1icIs2l/8FCB4e
iJonpQq9I4YmlT8vgt9NQljLKK61xBqTK6iTP3uE3UeND5KeSafUMdwX2vVhJ8CNsScCABLf1XPk
5elv1cYeFZKdOwLXkcAf3xB/ejzvjRUdVIVWM6rdhPdc1+917VrMu5oNcbMGpjPF02s7Io/ysBJR
FUGGwVpqq1YaRU1Uc27Vh8nPg+Q+c1tL8n8MUBMKcE5UOlPIxY7EAuKYkqHWzCw2kkdFE6Bgr66X
+VGEG/x8SVKaysVMOPeIwXRZRWuI9N7YD49XfYFY4c1o2+SI9QiK4USqT5Yl5HM2x2HZRpZ6nuzA
QSt6zsvwmLeb1fMs8Y8ZQkftBZoJanZnNqTlE8ltOCb0nTDV3tr4lRXwe8+KwgkaW33xFuR+rSf1
a7rbOaKjAu3bh3yo0SclkNodqVcGOmAu569EDMeiwfl35BgK3v+9InIkGZ1W2l91a9ZsaunLlmOd
VxERmeM7/dTwgA11a7rmjCFTXDpCXI8ipqFYM9sp7WOiNwAMiGwURqdNeo6xNSJ29veYdVCTUpiq
aLESgjVETXHWjMm7qCnCNl2xEf1ujkRtrOfKfMSCweDBKK/MS1e8M0sZMfEeWyKv+ZiBZ6/YdpQb
2rNUhExhRS0OVEzdcNr/Yv6i69NzLQMzk8l4J9kr6MpH++iRHOKHt4K7eozcts2fam5xAWXyx7EM
zvelARlk0P+dgomBNgnO84n5w6Z07giTB3psOWddeYwM5b1kfPqURF3jjimKqt9qjfwrU2ynFxfs
w5oSBYL9CHuv3u7BGXtgcoFfy3u+ZbtfdzQVowPaooehyo/kSiBU2V+PixnhOuAJTNHnZQEkhMEX
IfSQAMMJG6kLdWfJy+aaW4TVK4W7XIRfCN9KmCuaVdd+Qyrr1fWFOFThUg6gBrfiI+5/rbug1J7E
H2LdDxxr+olgKN2ugSINxabARFdkZ89ezR2W0zjYGUTnwSc4Bx+lIfOkv2TnSR3E42IDWI5JWRGH
exEvlDYJUCAmLVPxPEslhtUo1lDrGIXrQboaTSKgqezGvZtmnDdJ3BztBJz/XMGKY9G4muVVJ0Ip
7sTnKFRH3u13Tfmufjjs2pmPP9cgv7mMbjJvA4X/IhA8BNQqG4G2jSi2GQW20pR1rFI2v9EwH49G
/SYJNJLPAajQEVSoQg5Ptr7+PA+TBYvTAA5pp+J7B0MTRThv9yH1Wj1vWKStUEhpfgMh122g7yTs
eGe438YW6G4YhXV8nGswdewipsb63WIb2946FQsKJg8mXY9CYFQiFr4XGrp3ADykPkzZPeQbmfjF
mSkD1MLGCuDNKeXG0d1h70GoJTlc2c9lgXwpY/oFLQ9p9RQWNn3Kk2VIYm7PNxoZDlSMXuhYGNPS
N2jSh0tDUknO1wEGQG15v7tCOWORSnAtHIHfJCDJLxBX2ThZ+8dRYlSX4Jlsp9qmzhnEVVba8pcv
5sm+MCrPEz1wOyk4kVKdQNrD63kiC85kisfNsG4HEc6TVU+Udggfb7Q8sNRWgZzdhv6MBXuxaUAp
CI88QRIzEPGhNPJkczO9VqE1Rw7Jl6OKUmkw6QYynQyvb0uhF0lKn/OVKwky9cXOQCmvJ81BZI9K
bzSHB5Qr89nP0obt8oBSe5htHWn8VgTIhd06uAvaSE2mYuE1BK45bOyl89cMUrH0396yhB5Kqg36
ZCuoSUcFMxp4dSP5ZQfRT5YZdCsN5nCdr2emOZ8YEVw4s2Q5AdsZ1lOJCob9EO0Wgfw/fqOdRvcW
v+dYjmVfuBD5pKoCqws+jeiTUdLbU0DU/44gFuI5mJIxYl9NxaBFIb0rlTMWTcuSmvC4+8JJ7Hv5
mjJ9+1DmCEf3mb4zzDdFmhutnoUryoVl40XusbShII1XCx12rWTg2UYo2vfodO4ZBE8cHXUHsvTs
LipogTePCps14OTZbfuSMFhqujcu24KXbzC4r1tS1xDyIKJ4Yueog5B2f0J0T9i1hEZTsSlIjHYF
iraYyyMz8wwZ7QzoAYQE5ZgGdArj+hdSoPbIqMDibjntcTb3uRdlF/nb36NgIKYK71ygjhVITD1L
5BBSNpAuP0wImpBP8CL5dW2GncV69NxVIJPBQ7IznEygxpUqaBg7zvoqOEULfINTIImt29ClmUmT
gdPhlEWRpeWQgD5Qzxyj/tZDFVg9f2Mh5X5VpRVAvSOhizMBovLFX1IS6F0tgfMk1UylGvj2FXho
E1hAFDPRi/G/Hl9b1Ho5rIwD5nW/ozxw+MqDE8ojZWNUrU7fD6VCljUFATPrWdpLSLzCXcKw9wXJ
u7fg5HJ3ef3nC4tZSAGxAI/24MP9ex2TunFiwjzQyzUG6Cro9HSfNbNbbITIOvhM8pUnL6r2nPC+
O2AeAdR8kAwIys0UKpyMSgkTrstPI+ebLVUD+0P12azDGe/f9yXtJvgDTemL1q+YIK6YZlRg3Y1S
F7w73skG+L0JvE23b8QEYjpbqTGHKAoSt/uDxVo6wS1iOE8X2YEchvG6A+cEQgCOjH0K7UnI6nkU
Or/hjbRH8yKujVkgwf0gKSZhT1wixau0OrBSvJDlv3Vt8xLFpNyYXMMSR9+7QFZHjMUHS+owV981
eYnj5nLTT1tuLhFQwQcEIHbInuk4YPrmTEMujY4BlBxbGcQ2N9zVzI4LUV2ahRwBs+umarmAWnoC
moOWDJ7ZN4e18ImsHsGoTqkjHeCiTz5uSidO8Ty5EdxEpbDw+KmBfKdxj+eMe2+JV0s7avDu6L7n
+YV4vo3K1EoZULvw+TLBfo7SlOFlZvgOL3+Smk1ESuQHyscZSc600Cnd0ZV6BphnwnLDZER2SMpR
lJ7tx/4DnxOE6p83nZG+gOSEUNyZ/dnOwgp5e7ADwEt62FwHrJeQOleaKceJeAYx95DTyLHStJSK
nTk1CsxAEzvsVfpEyr2g0BRL4D2pKLBw6eJxLj+vkjteVDM81iOZ8WWO4yIZfMU8oSd99Q8ZAqF5
4A7QbA04jvCXv49PlfkfNqXRZd85AaFDd1feYUj2Hl5RyP0cHxwgzwfJgaGIEx6vXAEBGgnymB8h
r1OjKNZqAa0I6YBgK9/XLcmVgnoPLSitc2HZxYtHOmwRqCAaHNm1vp2hp7GsSsO4luB1abQH6iZY
59gnzPt8s/be6EmvEyXoHgzWg6eceXRPjjF8Wk5+cPeDfsvg/Zw8CceuGLLbTDEo5yXLy/L1MalB
gcaej2V6EC2RdW/7N2Ae7LOusxJv1L2F+CEY7g/O0aQAx3mFedjcn2XuFYolJmp+31oxi2cFcfjH
oH3w8NWkN/hKRTW5iMZKkpQNzHcZv5zOeV2OLvIbHqxcPoJMGTYI1hH8/BdVLjJrXQA8vYTJnvTt
hHFrQIvQfVheVW4e08Co3BXsrs/63N5y6cwnMusg/IsIuzirVEh8oMw3yYdUKUjjJral+VJdctwR
s+Uzuij7+imVSwFLrKSa214XJsbALTCov1hI+DsceLxszXF98I4Xt1BQAEqdYJibcwVAfxAdhmvy
08VudO5JgFUgyrHcAxbBy1OBqXhvLUlVQlgpxhhY8AFdiY5j6cRnBm+6NyQ4SbeMsXgZA3HYJyoZ
VBuAb5mbizyYycQADS0zlyLTNDzayFK/0Xzx598KZZa6/Zrwh7xzefZCwtFKbzKTJZJEgVUl9F03
ndQ+cLC7xnu0AAk+SRqfx4VYzImlLJU5RZH+eyyoDc8sUndkDNAcVlCZBJL6AZinxS0QmoGwy4Lp
PGnmP0yZBdX+SIM/2dl/hqG+WZEidOjbqjI9g8qG//aGfNQ0fescJeVEOdakxh2y8uxQwUsJAjXV
uYuebI87+2+eV+QD35WjWXCz9LiUc8byE0X81IWi1n7hBpiEDzpQ32wrMMcrycUjGEq0pt/c3FO8
SB7q64RIYNQY+S9+eIytPqRzbLNrTumHTkk2j59yPvL4Rx6kLGBOqThpvb9k8E4aPl/U1hnNA1z7
13C6LIw3cyCkRg54QuGGJJJH3l2dH1uUbX1jMLxoaHhiOK7PGH09sW0ZTfHDiUTwVQJz4ZOJ192e
oWO5DEOXnPccZvbe2a54Pzss0j4nGJR7W7wmoKOm1VtJ6Elf2e3fBL1ATe8oygCXKFEaa6iHN48h
jVVJ34xCKCWIjBX/4fe5ECcUt0ZKv17lu+3xXSb1S/Hxk2sHheIrkISOTBPeauEvAXMlHB1be5F6
kRejuU+bh/agJ9p8ZCRDMMkGHWvJKp+37riV2JFEkCogu15JJPUeIt89W4p8nrFJxB6lGOi3ryuE
JphF7vOJAIA1jfE56ZSLbXzEBVA1pPOxIAPSkfJgIiUeHOvGZ/7DZFmBf7MhaRukgz1fVN+Eh2+N
js5sieZQY72keyWpGSfzCLdK7xSCLwhMuUCjK1l4Zp2t69f+VhezUv1UtHlN0Y6YBOC5ntI5fRrs
/ix8CiXg12ju3T13p8734dj3oZJ0j4fQKZ9dCUPXN6UgcruMWy8Puvhsb+gpoubQG3YaIbumvuXF
wBR6K6Ff8JCS405msUE1ncGL03gzCZ6Pvi6RwNuFljCAjDtDa+BBeDSDQLeeERgSosyuUvw6StLq
CAhjcbyN6hhzeR9rH2GH//LTmbxc2laAyL3PbjU0n4xJmYBQ/wgmucS1TLmuEQD69ZAMjj3IEN/M
ZLWXB4+V43HdhfX6MMZzX09o4JOdJ3oIvYQ0Gm/0ZLpQPxFhLMnNjWADR16/SQT0EJ1qx/4/HIyK
kZBgQwOhUvmvqvZu0dArZknQhZx6Ypm+pQvk0Ra/ctLhfmP0FNexN5zAyuEu0lyYraNrQUKIwF2w
zolJRmYKQfv4esRpVTwBNMZ1tD0rZmccHNw1tbUcnmIAyo1FnZOGQMlKcMMdGjQ2G/KPddVwAkpV
GsB60zTOrS4x/Kvf3Uz1aiblDRj1xM2bYzQ9BRMAy8xpax76+ymP6jYCfaL3ksftzJMwuKKrc3Va
apoHebJpCDsn9OfFt2mWAFX15bwOhPrwHR64w4NYyt870Pr5gz0QpybCNkkjHnu/hUKdZet8SGsN
neOI3pcs7Pf6qQ90LZopzjbHay+CMxWNLg0tAfUj8KJobg6+WWQTK7WBLpV8QzzOUoyYDP6Yohhi
zkm8vMX6qS1toZDwS6HzGcR7e4zKt/iHPSeKpQhxU1pF1D+1mIQA1pDXVbp4zB7+Xjwx0F4bscPH
NKzYyMhzBM7uk4GTMTs+K2BrGlxxPIXjb8lA8akqmcA520yKo33N5HoWBzUmKvwuYUlG9TkvCY1p
Kb+oS8bg0OJlAd068AdwlR06V3jmcXWU7IuP5GM7L/G41iCJO2+z59TPMbOYLbSvEVeH0xMrW9k9
we93GeHRnPbJDec2P743vAK7MJHQDTkFbmVHb1AdZ5g4rvOV5PeUDeLoK0RBDChYvg/drj/NaDDa
CH8hL0m3o4mli/+W1Q1om+JUYLWpvCNrCdIO6T9kj2iRfc0s9HaGb9ljQXV18Spx7ueE/zW6TEdW
JHoa4yTd8Ve6mRTWPjRReKTE+w4TiDFba6vBntUcItBtuLWXshW2/Wt7oKEBz384VI8R7QX7qPYE
7WmBAPI3JkXpHwDu3nceamwsQnpVWS+yv4xWXFRDBQobl860KwM91bEDEjtGoQImnClYJs6Vd0lc
CUrK+QWqmtEVMwdQCzaSR0oJNF0CvdBSdJHCR+Na5RTTb890ddV4AuQYubZZyHQxWdbMa916gDDd
sKqDWSmYcmXWOpXIylUmFwGji+10C+ZMhpXZbTqWjgdrYA0/0Mg8I4OAN1VEFaGIujLnKML95OkD
7NT+TftZ/uSqXCmePxwlSrO7CaLm6FDuAXUE9bK0B3KTkIBsApH9257UXA931REK08N7tPQPtlgL
kL40fii5uoJERy+7h0djzEJZ4pfuXjZOeAMRx+wmZnsRQW7EGS7tg3YxQqQVp9HMfTjRYhlRIPgJ
w4e1IN+qeXHN0G1tHjUAKVBYUrAzkz8cPJ+UeqyegnAxrIuX3YJ0XZhZ0VOJuMpHO7uYnK5m22gk
uBGBGK3JoerdfnUaMUO1wMtLYAByD8GijyVoWM5gWRbWz+1pS6TzXYIYamVXrB8FpxdrmoUN4xgu
bUlp4Isr/F/UWN7POFSwZSO5ZOjS+9OKQGun967WFt4znlmbv+8c54ZgC81RYukAaWCP+S9hWObB
peVmC3zfoFQ2lME5GOWictc7rKLxSorNfG9SqDB8OCdH/Bvo1bnRGEEoiVJsVhOXIHjIdOAejAkl
02Hw8VtVGQsaNZGdEc/EBgafoiOeAOLVnozzN9TL4lkZEpJ0uW0zQfyvLruvI6Y+X2ga8KXDfpfi
fkrkk7z4Jq8g40CwnJsaXo30frs3JkPlPlAfl7oPFPBvU/s7q2azc2ddczsUDXEh0tMWH5Nyavhu
csQk0Os1oJAXe2mB+oa5BTfkcgQJodMWTW4iRkxnkiK389HVrKX/uWTzSNcHhjj6KZfV4iBzDcNC
sewN2QzR0Xryjevu7LS/qWpRP6m4YHTrLxkTHh8ZE2mL8CIMZZPPYn1lZVSHWvQ3z76yc5VX8d6d
qxBfJ5BsnnP7QVkHnVSfvMfOvoHzClE+PP8cTdTvRujGHBFHcya0q8gYZf4txrdSJ8AzwprQx/jM
L25FgGk3QpaIprs+Vj10mshMN9KkYbqKnTdv8wSuk1nm358dCpPcTSg709l3iah4P9ydgNGnYiIl
OvpkNdqQSdiz0mAvvzeH9y1Cbhx78h+AVia+Ypmzjtd6yC2+0vusGM36hDKHgSHZ26OTNRSNf7Kr
WnYHmo6cdLvS2dF0mhrYbi6OA4XePmFCVRWXnSgjJjdBt4jJ5guIkoHemY9LgDgFDoQFJmEwwgoi
WaecQj7rpGmZf3mB4CgLFKu0IhyASMLOgYrHg18i+R0B99a8NWWl9O/J8G9GluoANuQeoIdn3Rhm
8KnYHIupfWHX6n+mYN2t5r0h9quDgGvex7HjJfRyCWi9J09owls3cAPiZBKjNfy2izVu5BHZPDpS
MWO7NrNBVZSpUHmKXaSUq842WcxDGP8918AD/GPYo1hwNq2zdYqk4cgNCz98auFJc763xiSeeobU
GoxXXHINTJKOLaUItZ7uM+yAj1nTmhQiHV2wO/9cUa55Ps16MNg89kvbSCmIiYZ0NE4I2VLVVgoW
SKJ+0loSN2gx/K4xos96d+Eqiv/JqVhvB9cn+xpfjSyBvdyvn9BQy0JMsdizqyiFppmpG1A65XfO
8r67blLUEDOHrzRddXvVus6/V2cVFCGr5ZFsBVkogLzQzioGwy4t2Qb6OS7MhutidOtA+geLnTM5
M2J3SGWGlAMx26+5bYdNmydUJNeHNsSsDBaA10qKWWYgekKM0zuVMe6J2565NGHUAB/ala5EQ483
7lapl3TqiNy+YkxQVBPvxRXHv7x3fw7HeHvEabPsNuownP6EK2JOrOWBVnCT+kZL+WKTK0vvwuYq
rBBzYJNLxs9ovDw76QT1zb7UFTPrfiNszpvAtkG6DVYDytqXZdzXKnAbW7DNBDrH7mRx6AlAUJS3
BN3569nixT5wgnsDvAN0bCRnJkFScTEOAkI5gbJzHVriCr0T0JRN+7SoFC+lDxZSIY3s9e41V8pZ
KZOd48gCChhkGmDgiZ+QYXDrXFJ3fZ5O52aXFf9Vju/3K8zfhI1QwwNTZbU1DJPOvR/4elUpeTT9
0feEj9n0ehr9k1UUCE19Y5nUu3eCCPy5FGSgiLSGOmGfCBg5WI+M4rcGLyy0HiHSqePbWGvzkoWW
GOPQ8bnm2O/1BOJQAOd9AGu47fvPbNJ4CWaaWwTjWe6NLHwu0SuNo5ZeCS1pqul+H0rAdk+H8YLM
WGNBbqKS0eFG3hN5ls2fyU6sThHxZGuI7M3Yb7iOcD4yl0vooVhm1Cq0Y3VI9SDfoIhsQx3XyvVo
W2gB5KKOuba7Az9jBUT9scD/tQ59WC9+SqJXQzoLZ+P2KH5Bkt3dujaPgkA8wJnfDlMC6wJtARTA
l0vBr9mPpmARbQt7IzKxyfY6DOUlgu/L/MGpLyRcM81dgxrcgsZdv8Ff4B45iThDHiLOxTdPHWJD
oXUAPyHDPMlQB/aYpsWN+DAilo7dNqWrzVxwhSqovftW61eYp3Md+dBTJd03wkzo12jhGdJxFjqg
rWR7PAJ+gTuvFwEOT2JTzmQ5K+MCS8SmcUURlmtcI5RaMDpXWifraNiY/bgkQX1GqklUMeohThfe
dGnd+DdrjZPsiryDZx/3bi0DIwUIC9RJaSbwzLZpbzajZwwrRLppwpDCKut7K3SWDCPKXX48pLvw
ECD29/bZKM24mwrtKupIpxwbz9//xEL2foJRLrgY61En+aYq+gruw6lEJjCunh8m71aJzFV+J3Py
I7wzG/GJiWlSq8b71axB+tvYaABSiZoiSIlXLN0deXwqmtDbImPT4bpFZHLxXB02ggCupuRAI1e8
j8CxRpS02Y1mEKwxhyVNN3v2W41aw1jGKSKijX/sjRyX4XbQ728AFcrfPPXD3nR8H3aoRJkLDupY
6mRrqr7jkilPBg1HLYq8sylYYr6rEkv3+rkh4/LQzOGK6aMLa8lXMGadzIvZcTgmebcUOiD0EY/a
Ma3piL23jV+zdbzxympPttA8B0rJzIYoz+gX5gzQu82zU5VZGARzgjZ4EUvJR3I6QdHe1JZU11EW
8q/g5iQLSaXUDBO0RS8GHTu15W0DoWR4pc9+GncnKhw427LTIud8Vt4glKcfK6aEyCCAlw4Le/mJ
TexH5u0jcjbBpGCXA/FPJL7aYq8dLw4Ib0Gy97qGVh2K5fnQT+SOe1TCkiikNOetDZpBh6nQJWtM
NfuI0a75TrMSiMnv/pGaYJWbJULVBSKUJUGnNVOeG/JLt53pMeOWd64Sfxy3+H+R892dCo0bIk1o
Y4kd9gZz2Wq1xcsDFpbzYcPd+n3f6/TXVgDklk8MO5410YGesT2czjIeAJYk4iUVTiPJ+L8QC142
DUAil8T5gzbT5s2g8XhTEJJIMZJMXUd0N0xtOQbj06NqNXkbBE/Du1eTN9+MOvk0+oTgwS5kE/rK
Ob4GenDgnNMXrR9Q0tKxrooLqSEA+BrPM0LobzNbNRj1fj3lIj1Lu8bLU6TXxS8TC4Jw9nYHQoe6
0PXHKfEIK3It2GJtGhzvaeqZseWNBGtgwWrzfZOyi393Q7uS9y58BzRm262zY5XXgOQN6fjf6Vhq
vMmxr75dWV2mzEwwEUPLAwvOd+7K0r/u8sD3QC3NAAKobNgyuZz4m+zVf3kkMbuagK7crJ8s8lTT
SQuUfqCG2+xjkVwAq1+4q/5ddmRCuQfQIESe0AJ221HhdGUXy2oMphNDakhtsBRWoVguf1jWtVOf
Mk+Wm274lbKUlBdeYj/Fa13+I8NqHxr+TiSs492UyC/FUiC5HC/PdLg4nbLq7di/kBiOSklbhqDq
oKSmh6Xt50BCsvs0+hfy1pzOmfQ+A1OADrOGtSY3Q0yU9Hgt2kA0D/q/kix/Ot26lU5IYxCXfJZ/
iZhBkvf5lvbI/uCXG0uKe9Wx1UQfdWQuOcSTCq98LgFJJyhJ3+Tstja/Ijp4T9LznA2ZfR5lCD7C
rJHJjKMkPegYhqfXjbciR7JS2LFs/vWL+ZZR/cfWdZF4exPbK6PMk86fgoTcJZ6JiJi+rM7gphy8
jZKo04NE/g/UXyL+Hwy+XR+zdzykbuxCpRrJD6rkFBxuaYpRyhrh/6X/wGPRSibqYBom/mAOLVrx
cdeFTNhhUzT5BMnnhzeu3Lz+bhqMlbrpcCQS6497CIv+1qguC9Wf5i0mPwExKxF8VYYjcqMSPzEo
6KCLcMPB1oXnlHiww0HoPxyUtPvRXfV1bidhEp9a6CoH1tlLwx303g2l7/qLCMyJbL+HCwtXhV2q
DMlxWPgozaSsUZgEY0K4jClPpmbNvxJul8tY+dPxkeIpISkUzG1XwMXf66X3ai6NGReLAUz7snTp
/ixO6gvELI3ZzoqBsKALiKv5DZWl82B5jHZYyU8WaI7E82Y7G+dZX8cwiFPdZkYwcHBs+d52ovxG
ARiCNKVCfrZyDP/RtVYvyxVpX1V2t9WajyINhPmevT8aNOUG45DE4aWg65LDFvrgRszj70HG+FPu
eoL5kgQ+mdpL3EqkIRzJJt+1bvsgdd+/R/hN+w5YmWYl0ebYNr60eXpAFtwS2wiviDK61hM+viOh
/jmJuBGwT1lLiIImkx2+9PQGqwYqL+ZTQ/1o4kuseIfpRsB9iPnJqOL0jtA5vgaK+XCU5koJeJ0G
ABnFlZZIxaYs+fDiVDu09OfxW8h1uJ3IRwvz94+WJjEZ6nWUvsw0JthzHKY09CcHBeJzqgBTOd2O
oZIhOuJCkOIuugLyR9cHtpkR3QB5K77GYQOui0KEr2GUwBK1Z6FxclKFFu+GSqcKkBI4XIEA03XK
tSUZbCGXP1+aKd0nANrSu8zRy5oMTdqn50P3mzalzTYc6KUyLK1ohVvX+5O9WP6pJ9+gltW0iWeE
B2zeIVtaGznDUdn4XNXTUH0AyTRsyycAoTpRvqSggznP9NFgZPH/s2K+bwPS62sSyfrT1K7CzRnL
Hp6ku5tslNqEC1hpF6kOtuksWXL1os++2WVmb+GRYDDWEK9SD6sjR3qE6idGsQpgRTikv3V3lHGv
VkmQKJNKoMDnmp+rkBGGU8Wrbzim6TMLXFUbr6UweW1hjNwEmVfvxmzb2HW0mdI6KegxH219o6ps
+WqidhzroDAUa/q8ThwKqb8yK0sT3ExwbSWOd+hNPj+BTD4A/y+R33uo9gL3o7Nfwqr8ZcnPSReU
XDPEZUSuCrbOwu4DEdNqn5dEOOQQnjp3nY5DQG52pJpQOxUKL4zZs6a64c9EHUm3gylbv7aorho7
xHdy5aybtwJRtnh27HbjL87rXUpQlLqlRimgdMjjgkPsIcEzfoN2B1wIFPPjt+Ahbo58BcFB2XXy
0wV95h2zBYgJl4F6Cl1nCHhN7sYHk74WC3s0KC/AppGiAKxymYxEahy/ay/bseAP+GNYkkxkHtNz
4Yo3vUxJVFQMbC0epHEG4nw1w8z2yHi8nF1mODxA2FJ3H2sjW0Al1CIAbefaY0mp1M26u3uRY1kp
ZRwCoQyC/wSc1OD7PmqxtKA+eDSkSXjRMYGCJw/vrF1t+MwLWt6Sv68Iqn5IgpQMz8aanJ0qlYay
SeeVO49/qo6ZuKiinYo7qhE1nHxb2fx4tFilhOZUX9h3P9PKj1KwMrnlKirYU3DUhSgyreYdJq4w
FlBI/r9p91hPq7h/kV7V6LLJoXGvBjEcUbWmtEynLzHlBbygPzcUsed61ocYCDM+B3yKuisAcIzQ
QEYNJ1Bf+Lceo3AEO3FhmUfWrAnsvsde2keWjaDyijC2LC/2J5n7C7bfaT04rCfPQxRe4WmaG4DY
gTeHtXSCedgjaSvyJoJhfMZdoRXIvX3ePlpu6U08GQhls+tUFdU3lAoMmrkS/FuSglpFOO+eryDd
m/zVOchdAoTc5D7rwEqr3GO97Dsuax8LB/aOnBXijOElF1A82lXa30xZny1Atn/cQAfJi6b6FAmk
/RjqaQSOffbS8SFVg4elKgo9BMrCEfAkjxryjdENr/RKU1ogCi0CjDGDEIUFb9q2U+jFUp+JwqkZ
cdFsdIryIMxuqIKaG/8Q8MvuUSWQUYs7jNW+RcxP63WoDW1KzvcOf0Ag5ClS/pCvbwmQRTTzvSzG
UxN6beDXHBP6FkiP2Sln8NvdGzzKyiBcLGxUXqxZdUVLxp7/kL6kgF6e7QlN1KpRy+jmkr+aNX9l
wGJZLlnn3+19WaR+bHmMSy8BkzOFWKuHjIMk5sb6SrStcQscGq8uW+VzuhQ1/5Eop/nQ4O56e6A8
OEDlOwDv0YzeBpBCLZz3JJesMDPMHj7JHNMxS9dDS7fyFy/a8TjkCXaY2LIAGs/TZ99fILttHick
qPlaAQeD5C9Kc6cSFARk5tHng765hjwNdfzgfW6+x3jnxqsqmndYI5qDWagvccEYT5Ct+mUb8C2j
JXprIq9ZKPXtLyH8JdCvqGyVgyL98glu/Wo68lLXgcISYnUz5bNV6/DmhhImWx+eSEZw9MtJt4Sg
qKP3RhKnj2DN0GDkjMGoFp02t/mJqeSKQYSN2AFhGPdmQDc81elAZMf8BoHJQosfNNXPmszrmxmy
FI0AIEptUe9US3hm7wNzQ/DV1bMQw/TJ94mO/tBujXrgxZ7be6HjxOFjscecMzr5qB9FdadScJu5
8J79kWpK28Ich+WpVWXFXNImChIWjvE/NQG9ADiMowOUkFMyGzp4wc9pV/v7ZWCt3dQS9u73H2Sn
9mtq6eoQ3T4sPLpWIzR3sCoUFJO0mMbj8VHOmXCvTmnsbMVZ7FnfPcUeq9YiIJBMT8UA8xjwucbm
4e/m6xIlmnlIV9d5v7TdNpE4arvH6V/lhcnDdI9tcRvQ9n6TOA/5DRxstO7603KCXEU/0+OSLXCp
kOWRVsFHJEA33sA8evwfv1L1/0ZfB/VK3ZNkHS1Ff58OKMmTf2KCRSfw658v3r0heyxyUsUZaEWO
X1q7Vnq6qTip90SNvwk+zGZTeyse9Gi7GxlqGLUjSEErSUcRpqXy3WllqY7D6qTETQFANLta5TJH
lZtKotomWVHO8c8Q2m8JtrZ/8ZD/k2ED1i59tT4xUbqwRSk5yC1mkPyUjyL75gk1hTtGf7wNUX8Y
BxyXkXUQkJhNBsVxhKOFBiNa+8tQkxsoBmIEchEilCCq+qZt3dyhg9eJtkHLx1yRl3RaWVEFDwXv
KHZGabSfn2V2AZ3jXPW9AYG+cNUSqdayQCb7pDmunx0Iu89d0oxUdPlr4DRg4q4bxZfkYiZ3Dh7a
sBN2P0GUw7xqJgmEswFWTNykgHmHJ3cZcEUppu787iomkk0SN9Qn7kKetJxxnZnEZHxnd+F33LtC
keRWGi/s4fr0iqq2+Q1pPIiRTmmSjHDtUezp0aamTYeU9/+aKw70X8fI7Ar6Oe7TcaYP9nektAeG
VH6oOZ+FF2ioH6se5m228t5DjkwjHvMy/OLj0C0QAGhK6WmwjLZ1JQ6b3/hUe2tVwldmxlOElgW/
imjnBqzH83gXVMSn8A4FLio5hHjIGYZLJq/ZjUKEj053/Ulie1yoCv8oTQlcHrLqsXoVS65nHiJR
mcSSZBZ79+RacZUTVpHi2hl7QjZYObHH7WJlRC8ut2pEoH4azA+I3KKAL8VF1Ev0YyTB95g0q7JA
BYiksgvBx9IiLelSQxv/LpQmrMYWh8KI88FIuaVJ9jedPRm4f75p7qi7UDDbuL5OZkVjQ1Y67hti
q2E3sJE58ncoXyVZZBEfOp2Vj2h7PYwsvfItXJ1Ny4DJBskjCkEiuajz6NkTUjNZM6F3lpCEwXYt
17ROyAmntnLwybhLGthSTw40WdneGATb1WvGYL2dha8YbD2fOqaacQDdc20v3B0ZIQar3L9KBGoP
y4s/VLppeuMQlncnhFrR+tixWJ0yLi04f0OpaCiITXd7KJ3nsqNPTZHtIyvc018LokPNU2jRXwou
rs2n0fze4sKuyOUD1Grl3U9yevZ2rGfRlRDD4fbssKlXSHjD5zcA8J7hwLYGwvcJUPSWDPdqSLlS
E4aYry+HRTEBaKS2qDduirfgeVn9FTH007YONaRv2KdRUUhR7STuFYjkwgxCGLLY5SOEkAqxX8JF
W+bH5kGH7mbWEnKZnQ/o7aoA14XdJcwQ3jwhODb+k3a8q3d4tYy3GDvHzlETvPNYw3Iz+45rWcCv
5tn6rClK4mTSETjuxxqffC3rGo+pmtualvBm/VhI0uRrKEdkY5fOXjtzAcjTK3fCtDD0U02wHupS
gy+gKNtl317uFktIxNyz8IPgp+aKIQD2/nR3lv5L4jX7LqdpmLaoAUWBuoLY3B7V8tRX+qo3o+Tf
I13Mt4FavHhHsKihF0sx7Ryc/GTrHO4Uq3FQAyk4ko307tmpmXEu7EM/t5RvZrhBKHamSUgagBHd
e/w6pXEgWHQwy28HFEfmpgLD5gweB5UqKE1s/9/udRBWJiRXc3sLLcTga4pPhWnsumTt3rFhgYJa
KOCbm1/Cm50RMKxXQiaq6lonHX9szUV7/zlzfeM7U4vym+Bxtyt2YtffyDtr9OHSQnJgetkyNqSi
qW0SMC58ZRWETshXCQR2wxX4rktgXuzZQNcsS16nmWXp6RsC+okmev0iUfclbmEMTybfaxW4oJXZ
qkDGTwxyjF4b5NXz0EyujDXDiq8vcyllrZmcOpKAE+3iL3D/XjL9wto+BzgG/CAdye7N2Ot/10qJ
DkX9Hy0ucSrmqgkFcb6GQrvmCm1+AT5FVecnDnV37rvghkyzQ0M77rmh7JEY/NJaRXvj+0wWHiIe
X3jYbOCvm9bZYgJYzJKVzNSiuZ05QPj7wU5S/WNaHryhL87N4iKpSTo78KiwNRvSGS8NW0mOPprR
I6BrCljt+CJ0LlQarTSLlYZ/51fyPs6DglBPxDpdrHwF8X0e9dKJXkmnlUAdfrTfYwyx3KA6l6kZ
KBNEiRFpmsg/SRv2GLFBsA2kU74qfAkFN2QUL2gdqln97FXHzC3BCqzYuze4Y7JCTyuIxgN0RDFi
ze+unPi/MSQrRJbdRWsxenOk/NRh1GPXNlZdFHsb8Kx2q1RSdqD2U3VumhBvDz/KOmhcTy0Qi4r1
Q8SaVb5RZRNsHtHLg7S3CIRnzycEYBMjOJ0z2dwCuIaH842Wjf+15TIhEGUg4Qp9vaMT9XptufmX
3vf1/afw/Qu/bkHbH+1nJXu+pC1BpdiCMm3e9aoL6tsSZaqyhJim3AAGAVYn5Pqcj06G2bK3IcyK
XALY+ATtQqpdUa0JOVYTZbv16ip23Y2DsyV3/VTdyJBs3x/Q5o3a7Is2XpPHlmzPdLOEr4LAPA/U
IU/hO2OZTskHP/eSEMRYcF0cwtJbHRSqkbt2/bzmlY2xgc0zQU+JxGa6xny51qKKcBMPmLM/nSrt
Vi/50+fbgnf2YkSknl7Q4h/VHPD+tgaExxIGaXDTcKQhvYapIsgjViK68p7IhyqJdslD23AHhp1S
Udy1HzJoP2YdGCEI3gY8yepE3aitk/ZsB50y7k5TC6IjPuKLdwKEPTGk93SVRFerYdhW9SwABn4X
7zVkX8fSMtBEdAKY3nbVjE7jx7wVcz02WGTytG5IYzYtsP1Err6H1Q7jHCqjZo0DDDOs/6bWLuHR
aQ4JGFwMDQOCassxaggQ2lb26VuPXuQS3AF9mWuJZ7m0RBzFk/039AW8eiu5gZfeYua2YmcXEe0k
NeElOF3zY96fggD3AcHLWH1Wd1vM52VFqOmRwG9yZWheCnziheuzxZqf6qSCQwj/bFUqnz+63UjE
8eH5fwb+dhA4ONtLIrkOU6dwY0/SJEbNrd1spocOp1j818nghrEPQedz0MOu4PSg9Gcxc/EpLQOQ
omW7tlwcwRRX2kNeijOgAOmbrvBqkVpMPgszcjMzcjgqAuVhO12lpIPwvWQrxB7Tv2uxnhioU+n7
4rEGvNPKF0NFfkSASDYz1BN1EoUYzAp73HWNbpLzAhc1eZA/PR6Ln2iotgMA+sdFadfdlXo4qy9U
3ukUUr8/dPhUuahVeHl765BczUpHoOYTgIU6yrDCULhmxWvAutQbTjW5r3mHl3/C+E4B8x6tRzTN
Ve/evuPMIzVIWjd+z5+OFy9p5IG+zRwiXCl7EdRTWyb5Xl1wP/t/jqrnXXsYULPWaU+LSQXFTPyQ
ju3Qyl6OFYZnik6/tfEy79CKciIrMYTpDbTWuvxFew+Lz2h2x1lxzAi8wIchHoOiXRqDJxGlK550
kYlxsrl8yAgWfxrFcCjbgcRXTTa6WFKr+PmaIu5cfUwdSyeYEfjNe/xPevZYuVJf1YRkE02z+YvB
vJyYW7pQd7J5QBQqPeDxS6+sO7uU2iw2bbAxVCn3h1IsXvBO9mi7tZ4r03eVQnZ+m84dhqa3XwVd
zvGMZpXMa6U9ffeoS42cMmP/foZnEL1XyjRliczi49FkBJSbgfH/Ip1xTvY0z3Oq90bIv2EDmO6q
e1fqzXVj713b/813TJVj9uuhFAhTfREjsiPWrlXTymLtRb1EZg/RQ7CdjhxsBYeF81t3f30ePDvC
QXYjUc0P9/gckM/Ha6jj7tofK6kS8ReIh9vezMoJH6LEhI6o+5B4votYhK2nPftQO1cz/fsHPReh
QsBThLYQoC2Dv8Ydqs4IsT7QicNdQg93gctn3zCSu10coErIGFG6LnMbZgdr1C1rHE2pI50NFi7p
LXby4XWHZk5OjjVSZ1MKLHzJvAlNyc3GvmqR16ajAXeMLLP4BsG+I529eDvpsDsXcxcfASRvhkFM
bxH7ZiYOSO3y55kGWhy9IcfPYFVMWHjQF65LYK5TwqWduaSToYcrY2WT9UTsGR5YOuByXF2L+atU
8j43Fumm53kjsuAMQ6gDfLpX80+qWslF5HE4ZZFJqphizLUolI3HB3tMHJi7F9odMrgzKMOlbwsd
rkmqUnNtgQw02vdSsc5/9LX7yKCncB4fOjbr55/zxRx0QcfDmAMT2OLRooDiCJY3LBqX3P5uYVFd
kT/XTL6aHHwFj6l9Zo2yJTpAhERoMiZTZNOlyOrduWrZbWNq7pURz+Ea4bUocEZYPvKTYl5HHnEa
w91esb1D9+Bj/zFv1ogyKJhoFR99bX5mWp37Wrr6xDCFnL8wFjyNpcriyz3PBjxFR9ZRluNNcCe2
VQWRxDyRAQOU9VmanDY7Ei+RM7J6JLN0Zei+12ay6k3eL8P/Pv5hYCYE08jMJQcRLqcm4errSLx5
ZCB0ArmZEcxE7uETECkTvoYTG+UJugn01yphUcfSi+rxHREBz7URjztR9SgqQhPEEWb+DuHsFtd+
p/NbefZ4TpSm5SnnRcTbQn/Ep7lf7AkSKUIzw/FBZyJqF6df3Ga156IShv5rVvp1SG+kgKIxCKvi
uqb0pIszL8vg98Chq3iN7E4ap2cO7xKzbT5Pm8oJegkCd3lVW4lfsESZgoOIqt760lHyMzBxvrV1
J2f9sPDAtz263w3cVDzMEuKJaxUlfpBIw5Fhxj+kKvM4VlCQ7eiLvHV7YOm5Qf2716biKhr4oumd
1lM5AkMeIcZxE4mmICoqwOiY6Xt3468I9if0JzEoaR4dM7XZj8XtEulL67kRXnsq2LqIyjIAdfOF
k4UZ5gRW8y2Crf/bMp6qJxFUtoN6pINhtLBsj8GfthkIJOsZatcRB2NxL5nYD+5eDsxZwMd5yaFQ
2UHRlH38O5Kp0eSaD6zzIj9NxMNbH5CTfcsQq0LWDDwf3WWCa44iFMK/R/Q8oVuswk14uyR0gv6L
JwGIbqCRjpBEdeOg/yQlCwQEGVAZgpBt6RfHFYDohckUcmzjgwL3m0igB5HArfRs0O1javDbL75g
vRF7HFEd08mNoN5Wfk83+DsXf9D/dPcge11JjmbEWxnY4Uz951xiTD/CoOL3NaxpxuNui3cLcU+X
V4q4PGyj4zkJ7E3vSi98usdx91b4AMqMnaLf4z8cZs7lfvMcSN5+duv4YSj/q75V16QYf5BC+KA0
pShWMj9Wy42jnjkZFPvfvMhB8p3yJDYN8MFqZSaXSojNKwXbsuBcsY7iO1Oy1ZLFmIKMQifd+Qtl
K2Nnj0NEI+aq4EpHx6qi/Z1ol+oFo0nwp/jbWmIV3VhfLDBWmpCxieO5XgLdpNcM3URyt9kwnZBd
Xho4TS5Gz1Nmv4KUEjObfknmj2Sc2OBW89o/9Ts7nCujSA+BYI2wAo3RDaApnld3aLvVktccEd8f
uzrdSHpQVRRFSU4m+4Gza2xVXcyHypKaAzelWlHO6vk4k6c6UpEbjCp3kLNffTP+D/k/c6a4P0sA
uzFz0UVFBPkXjU8Fn2fPBed7UePVfNkOxS3VUBLVTJdTFYg9f5hVOL4tz/YeJyw8hDfftxx2Hsc+
Y5/2i/f+SZJja5UEkK+Fvhw7ZIh9LMueh+GxYLK/khiteUVx7sx2tsGRO1dpMvfet5Gp1wrOGTv3
qditI4Ku/QFE5g/cHym3gt0wJ3fzBwG17U9FsWu8kNARKWKj5tU/NgCKz/RBvzayYpvnSLrk1dkf
8frtVR9ikp/jqIT9zCCRezG5Ddcv3MK0xYCCI5Q+FDvqR2A5pxXZ5zYOLoW4bJK+SuMC60cMk9s6
/Ve/5pjQWHT78sTtaXzZ/bhHkCHbDwmE96PV/ZQE1aSYS+yPpbLN/11GP7+Tb5KQGLmoluvfMPhT
kTngEAtNu6IBvx54Apo9Awb2aM1/fYih0L0fYkjC/UhPYmPD6JvUU1LvagpRVB5cXd/Ax5AAmuDN
s/wTrxA6gBi9v/epj4sfpC2ZMQgM6LbZ2e86yw6SUuwTGkApHXoztF0+LOSaRN998Dzmqhz6jqx4
t+Fvu2Nqxl2AsyYhlWDpTWXYi/dZb3AiukYTltWVVm1sr3/MCGs/lL+/9t7Ot6lp8ujMPGTefDyQ
kDqjnGIDNziVDCvGNbx58hoUx8XLFJ3hS6fhh9C5ZvkiLZOoB7iJQ855+PNgWQ9spzEHRyYX4Rqa
aFY2MieJqJwV9f1yV70BfOTxtQttoXj4xS3BRXSaQxn2WyZCQ0IO8uaCMwm9cGJgABTW13h5DQYV
1ZzHWEmVPTzowuM+5qiIcU0zQ9s9BL+IhIon3Po4r/CAikNB/wtl1XpQSeg1b+RSCrTsqanBMhc4
kTvXOJ1DFnCV81JLqu0I47jffMnlOSAZN6omisZLqMfwhGcWdRI7srEMrHF0roNELi0+KzNcVia4
qVPCwtVWkgsZLjLBsVQiV1NUvGllyzyitjUTR7QBNWKiJLF9lFKNoOtBH68hDU5jV9AAJ/zVZsJL
zZnBHvQ6y/6R2LX9Yez104K/yUvVyX+X730nTITXUhHdLI58sMX3ahxLR0b2PZugUUQMtbFkyw0T
NFxts0hHA+wPsp7smvwWvKg5uXJoKqKZ9M61gcp9vTJks0lpJApWOC9bT0WUoauzs++5tMAnyz5S
wJsjhrVh5W6LIwYai3jTloFwXyci8JXiPl9QVLJmaiS0f32i01mM1r1cSLe7Y4K6PJAN+8SgNZOx
aUdrOjSlhQyDqgAFtWnLiUQeOyRnDglYCRhz3aSDTHnZ6WBkO4KaZT8BPxPYN4WRpHz77c8K7Kt/
Zb1cjhzYEure8eLLA7EROfdGBGSn8MziIvrGmx4qjmj/rH5+PhMwS3LTLQesNveKcBz7GxR7Z0wY
2GkeEA40M4PhO+msqUYm0CHKWGNAJzEMBYTYzGyg4HBqAmXiCq6rC82txSxKG4QWDoAvmnYsrt2O
4jOAQfOdicLdxiM22PZbwR+hXiDyWsXGCG5H2hesCxr1gm7v8E3782SJLAkwcDK+43+/Al0bNLGk
66mf7vuqJQ0pk5r741vmwGcyRAIaetr9BKF7+pSowdGloHaQSGbQOdDzQ7n95PfJC6En4z6ikL/g
/47wU6SLaq0Xf83aW1QjvJGbXSnfXiNbbqF5fpOzeHu28KToN5VTlPtCPEMSxs1cX0X2v2auoxES
IrteyC9lrkPWq9pyrav32El8iyM8ct0koYFWSutblEwU6MMei32lugsIKxzMz7vNB3ru+QVHRL4P
vK/+tAveaZgE7Ue0YXgXldd9I9XdJvalDBahC9ED+DlrkiAWb/dcNIRfRogJ7bfc7Y02g3Nq//4n
RflfXR9kv6tdHAr8Wz46QtJ5eG/G/MQmZBep8qtqJpp/l1Z32ifiRHV8UVDlf88u8e3WNxHfqji9
lfVqPyHNWbk1z6ZzdlwjatBpH6+sdq6jJNNiJbzcyvh7nD0NRFbObg+edNalv2yCyoqMGy1dpAZd
Txud1bE9ymgIqWezssVIfLaTSD3jN5wIR/SyiApRRW0HoZRHbKfQmPPfVntLDfs1O860zsHZGcHh
8t6scTdc1c+nr+4PIcsSQiNIPC4nmEdwukoGWyqON6AVuMWGq8frza8+Pq6sfZzoP8tCUC7EhySu
x4q+myHb0eBsxyWsBYoMFxeAMrx9S+KBJzi2YAxHzJAJnMoc51WRnGgsSsO7hi/m5zup4JDA38NJ
xxyPntHxzwY2/vKjSJK0/H1w1qgqvVYf9bSzIl0OPSf3iQKzBGYRrAwxWM4Z8NUlEyJhaW47gkz/
+lHhHRBmJzDYM1Rudtkdhl6PaOGF/ykM4UpEgpSiKHYkQO65BJn0PMQ5nEBHZsVcJuPEbrnGrgKl
DZs+saYD8lbds/W1wmt7XhVAXnI93axm/detn8Pm/2Jw6BlYvvLnkUruLOG11lhHBYvLIpTDj6sX
PsBmDWyvlCgXsX9DWBingcL8Q9vS409H4NlAsvXLjnLpaUzKbNGoVJDU39c1CEJAYsa7+MyvcDc2
sHZ/ZyEKT/1hluegXC9vCtsoYYBA8LCvocUxcVjVxq76w7gaFrjVP+aRABZDGNrTYWpe3hjV1+A8
jo0u+SmsjC1hCCg8Yc1PgbpE9FM5wL+2AHBQGkuGlmh9GbAHEDP74YUmULQ9Nk+V0mDeGal297dQ
mvLBL86+hqeJjcEfP2JL2FbdEygjazf2QJp21k+JQyDK+R0e7xnM0wHnPfpsro3yvedPUqYgP1u1
VxbS51akNUYu+gDtp6bCeIiE2PLzM6kqbVKB10Eb6mafWGqvZsmiEyBTph8fQXafQkoGy1U4lmDQ
VZuM0NoslHOiLIQdW7tUtnommjdItVFkR3oWmwo5H/ouiCUfeSpUdAjaJ9rdBOUhVujQ9WAU0CkS
d1GviS3Iq5BwSw9SuAXHylzcsMAxLVvGDDckU2u913lSS+ohQyS86b/z0HCkdBEKjxjxSRxNMP0X
Jz+2nFSIrDLv68w1zVTNQtiYxHrp9JtIy7IDjWh1DQ9wPEalVrdVlmpbUQ28ev5bxOp5TmauLnZJ
jojWtRdGuA7AlCcP6xde5tJ2WKQMbRi2Jn69YzcOSSWbqf1diX26Sl5Gsm0iryGmq9DsfES2UFn0
mAOePjC356zQjgyRLxBxmQuTwPLrnEEJfhAq7l59W3ss0HXoYyUd7raJ+FwIOmVjMgGfVcLvkkZC
3k4MGo+QG97zRF7Z17yfNzHH8mAdCeHwRsELn52hF/C60hL8aIM9UsfxUhn188Emxu45FG2pmo7n
ZbxdOlGwKHSfh9NG99w7W4rJE4rVFjlXQJi6fUFjrPr9Dyqjl9MuFgtRl7ob7Bogk8DEPd9bzyAL
O25RQAyUPe1vrDVfITq+qjKdvfmdTsdEznqN1BGjx913K/wai8ZI25mkGG44QzY1pBXMb9bpWMmw
ehhCKZThFMO9L8OXuXo9BP4XL1Avhe6QoKTexWE/wq2q2leIg/EMc31Gm5LzJy5nG9QCS9Zs7l5K
wd4iqYvlvAyWsF//H5UV3Xlf90l7iriy6HpncseECwbCjeBT37Mf9XWprvS15odNwYYRLXHzgkz1
StqJLEzIMh1mLus2rkE0YLAb8r73pUtRrzeJBosy3N5nXgYo5b5o0LZ3PiKYJgr0i1Df8wxQ94Pq
L7X7hYXY8lXnoDhvAGVafqJ6zPWW3t3WdT4V4oXulh08oljGbjgy0i9NSJDpnpGj6XCsa5tzvwCX
C3/eWtqnV0jNlHL6pd8KOvOGnnZo3cOrVx32o9zXqGjxarxJuoclYwy7UF88fwj1eqMzkUxj71FW
V4t+PRvODVJyny63LiReotgxYBGj60c7DNMcBoy5ldw/6S4WjmcqII+akhEgOC+3a5KPPKHGCit8
kYS6bLew2VOWM1H6aiKMVgt/feAsaURfWmiiqPB+r438uIkbu7a+eycc8exq1g30Gi2IIK0v0X2n
EbSFFbKdE/Ko2VMdR6ENmO4rACI21vN6jWQB5QfBrPfhQd3JlYqoGbNEtKriK+OR0LsL00BuUnAZ
qYiMGByd9aFW9lZtvo8yyG4M6P/L220i39R+xAQpYZb1oGZxAhnZtv1/IbZ7NScrjDP4z+6/etAa
MhYjFzUoYEuzeM9zk6RjQk7sXCV5/t+BOICFhjWRKq6QBbijyX2+f1DefFhleHIF1dwfUu03Bndq
CB+vdQoNVl/Ev6mFZOJEJ9IvSqPGRBh9EAErqxd3NsschYOOFDtftEYfezkGMkPDGx/otMYdPsRn
mPV8Pv1D4qOAdRdVBBM9EPZhVFujcB6GcRjUsj8VVZFzPS2Wgo8oKslfGas/Rd6Mp1sQdtgXJLCm
N3pu+mmhFamPHbtOV70P1nGY6cWTXREOnsUcEIfjAc2DganYmdI+90hk0czamyDtCVU+oXew8xXX
PeuCeblj0HDOIAiZKmuS6oHeA8bQrauoZttGZEZYZTBGTwtxkj+M+ASdrqIvZLtlXAllKb2b9tA4
zcANJssLTJUYtgQ7gUt+70xlUkt+s1pKK0rw616xlprRokec7DeDsok+D2RQmaZ3snPyWwGuHhRL
5HX5xWCecVfKVyY5WWxCRyXRe13s9UONzsfNtFfwhVrV9mwVFsPirzNhdjMMPXwvtQcJ0yog2sr8
Ypexuq36QtNyrxZrRSki7N+jdFaBiV0DUTGsZ+PN5N75u0Chz3XJFMlpOXfjE3Sr2ZN0Lys11O04
IyePgtX0+4lNmDbkxWQC7XwrY/ipfq4mn/AvkGDRECgWsOaHLnFahB77BFsMBiMax+Y513EyOc+m
mz8JB9pLP1D2hQQ4TKeNTGCZIsYUo0mRxVvg7zcsHdnGUYQD8P3JYK1yVBZ27ogJnwFyZWAi71Es
O0BfmXTO+kA+p27pw01GUM04LpVt7mudDTivwKx98z+mzo2gdVxcDe2ootLXk0fm8H2BpTzeqpYL
QE29PpxACAybFZ4ME/OzNUKyjc3EsgIs+2sTtwRpQbCn3ikF9gfsv60/87gKhbGUAVkdx0ZYLcpt
+OxCJDF4zjUzGxGj3JgE186Y7edF55hgAMqtUhcdwOSj7CaK9yc6IX/a6wCQ6vSgzwXkdxAockob
ZXt0FPsepHKJpy3JZAQ/4wwMFjXWqoGFKCYtVgyMRCpxeeab0AJ+8i9xNEHcNgNAw9w8MEDKNMxG
GZEUYLjh3oBrZ1ggslgdb1FhnJuyvGSHFyHTSTuyy9pYDBp2YchpmjW8o5aXmZKHJEuCXP3OCKr8
ejlq46Ct51VWzhrwdD3L8c8TCAC7K7vZqA/Mvfbp8Xchswt8YZNNxjMhtbFCmohtcSU+2X54q17Z
0/fp2yGY7cyyUIWkTBZubIK+IFnMEA34NsqQhoJwVd1QsfI3fC2EyE4Zx/04e6PwOIac6wIiAxTI
7ZBRc1zYoIxW/uso6stjBppNkOXMM1b0N8QstbTB0JT80BhFblKKyXRZlvNly8gNhj6VzvWr2otC
1iOVperUV1H3rGBfVq1Y75YcJz3eCV3bQ3Fya7O9QajnU2B7qJmSHlARr4YJGb+mMpwdvln/GYeu
+f+msVaxhT62gM/b8au4/yOxN2sfshwE201qEQxeXV6cvCMUNQQZwy3eFhD2umguw6bq4d6Pypdh
NbdfQJPGQNsiXnhOFCIma2CfHmV0G58UPw7GJo/G47VUWIM+h2FsvpHa/dc7Z82y0vT5mQw3GrLk
qWo8yT8f7L3h/pKZ1znzpeFgbSjHPNDgqdvQCKfjxH8kqnIsLUy9btefAC7RiUDeYekQJb6sWaw3
GOM+BtlqwLaJgPiufW79PbQ0ootwrbE0s/7dnFM8QCObyT1QPL87genRhnY91JBSYT+XPJrxbQH9
MUgaPYGtScvU/R4l4fTbOlCRCGFKYIz/xPCAo6z6ir40mIhL0bmbAf2xWCQwwm1rpAxcKJNAe4xF
c2NtUQ0RecaLtnzHcuGDHJE6ccIfXi+XVnxj6s4HUKeaO8j5RHgc3wMbW8kRd/7PL7C0rxbuvIkl
UuvM5ET03lykosPVKI6WAP5AlaBKONm50pyiapvEgedHYmslggEeLejA0MdMoeOY1A40ton1zfRR
IoC0DX4WrbZxZdcCL4v+6I8fLDzVQWPhDRQgskYzXg7BbRMagu34rCdTrxgod824dd4jmkr3NFE+
tw1dtDc/MvL0Lb0/NkHg0rWYxjSA0fzbW4e0ESLPak/3cb4X2/lXDeaWqfvzBgjY3grdMzlD7Eko
ZJnRTrvJfOv5BpUDqgx/ZjlPsXF2IWB3D3qUPTNwIPONfpK/9aaRfVOzd8qd5Xe0HlQOIla8BLbG
61EnwzjyHsgfIHCcm0BdnGiW3zUdDeHG0Nsu/hp0gmF0DUmIctMimxUPglt1pUTgoiExzRsregtM
dZLoI2IQJUeGDt6MuVk8DMUff4e5Cw9eA4YEn4RUkpX8B89ibFjsBHETPonzqNEnHt+SvlFKEpGW
LzSp26uZtRtMplurTUB3g3AOEfb10r6mMfICN7dMlhzi5Km0+X9f0AM2uG7sz/ligkFn2/dIp9px
I8OsFWQfEgj3E+LnFIWPK06RrI8W8RBVub8AderKDx30+S54wvdgJCgS9E6SCGl7fyeSsgTHJppv
1qogCHBiNqa0SezOESpY61xHtRkG6AmE+KG+dMpF8CQvzLoVuSfsIvgMlKSzsE9y0g0EPTULHP4P
PnkbdN3Qk/RHDW1FxVp7/Cq72Doe1a26GFABOco8kPr6lfaiK8DLDB1EQgTX/nd9KmN/KN+NDuFP
kBKBaykcHB/f7NY4AzmxePHXGt32yisMdfaovhMYmaHIzvlsEHEnj9zAgujnIkrsiA+Rj150JumY
rTdvgw/Laimxw+SGG/mTOJYFIVsdEMKrnUkE92/pulczz7UrOtrrAdF0lR/35LTb0NvUmgR44S5z
hS5PLw2zizWgLZWYL5LTMVdUtdY4nQbjCUYrwoTTVGcP0/3EaMD1zatgzV5NKw6sl57V6txJhXjT
MdVhv94sjfDA8ND4Ewr7KM7R+6QCHjoM5pQX2CjQItJojJ/WVjFdFxHdXrdt1NlSruD84hqD7xPr
7CQoWtXOuKyRdoxoNz83LGDvgnqjW3T4SoN/OcmTvp5Z+mPmEsCiZ7VImRZzAXjW2E6h6nK4KwM+
4goI4iCCUsXUFut8Danb4mrIHNWyYUOrx6uY0K7Fq8tha7dXpkj2Q0SQN01JVNiE/iVPfLUxpIt9
x0Lqqu8mZts20E4XDOA1wnYf684WtL9XLLRn2QmwhLc/vvAp9cbye3ajNAYJB9+QBVSlbgVXLfWg
auEV8BHe82rx6LaL26tCKs9netqA6YG75lnxgv2DLveMTsdfFl2++B/gaEL0MCrSqjFYwf+CQNjO
O6vqt7rW58Wnw0ZEGywVfIMBjZBSGmBsy3FH/nRYXHLhliXkCPixKYA+Pi195oQFkGE/KjM3zJu9
1/UaIRA5oHz77UI3QrURc4lWUEAP5Nx6t39Iw2Tor7+GIkJWrCsKUn5ffa/nRvC0WCZAYBctsRVi
RQPcSdGtQLdqUSGSCZVLIWIpluZgqKQUQ7y424S07VqC2zUMBkq04ajzkWbEUNe8Q6lRniv8dhmc
Hsrh1Bkrz46rRlwjiGl+1DBQyuwwTKCTpOJh5jlUAde9OQZDlXWvOW06DxBoM29vFTSCIYRkWxq+
kMDn9DZI8IKLBEhiJO9Cv2j3w7niI4sc/XZF07ZuoKtch+ias+4y8HYxXxPJc6D2U9guJqjcXZ6C
izUMFDDd2Yn5CrgD8GkDEyfG/BA14e9WFPHXGLoDt0Hg/eqUoa/HowNTo1i2+cpTkEZ8gEJFgpbz
NcnXrMX2kG3javwafygRQ9wIMz9aXcSXMkYN34BD7AQ1FoqQYQLsnwVQF7ZG5zpsBIUmKPKEtEll
VfjqxJ8sKeW4IzB+aql4Yp1/F/lzZNuQFQyHK8GlZi1V9pIDLuYJrzme/FyZmIYujCpXnPgAR1uk
4JFRhK1Lz+VIXwFb+Ioo1+AyNBigvUNZanP29J7S52w+szAy9Jdy3DYKu0M+i6ucCxD5GNzyih1o
mOXFSZzfsD0Ehw2jbIZGISnq9l9tT/fY+v+k6Yds61+MO5rLALDFFlt5JN0dCg+gaqmafbETxwd5
viPGaULeORGrvcOTgVCJL+8SYNIKhXjZ9oCRTWvxIWJlMeQcmDSMXePM82F5DYi/ynD4FINm/i59
j/URCFfO/rw5WBBQj1sgdIVw2bkS3jim1YoKTqtvmnHiNp8nT6J2cXLOuxIxnHaoQ3VZfjmXMcDL
VngAsk+A8JxLBUWZqlxlStvxpRZZWhb8pbv9lWg4vmIuPXlVnz31IXOTBFzY6x6YoiGUhuVZ9GOf
HMHhPbZIUWg9TpEtTXf4WWUEd6VIyf2XmGKs9OQCGb1UMQ5zyb1MeIa8UocnXZUmjxL9p+ALyR3h
XWcNGBac3pzqmWm6cP2gwCMTeu/GZYgcpIHCphCyVuMxsVpz5Lv4jq6X26A6j8q83YkO3ExdYQGw
ZyHwMVi2pk9DPjiFNOTnJi6N1uibXSANxB5GbVVlxoavW42kfHeZAQJ4kaRmn/PhifyPpeQ8yNHv
HJe9fmD+Jug5sD+DDHX97PiovYR/bz479AufVEUTb0BIi2FinYpckX5m+vbkSG4KVhXNVC+37ZCm
f5oiQYqpl1u4v/SWG1NLCbCeRdxja3DanhC5L2THIpcGs0wZveZ6NfrCEf7H5l7uFO929LDgQgjF
dTbK9tx8zboPVdNfb8aZ+uwhaErr2vkLJHTQYB7YMnJ51fiK8te85YlVfTK7BibIHBAC+ANfyv5K
jv7QmSXPTeUAWcQhzenPIka6+J+pLnzkriHy1ywqQ2XlebjYUx9TEVjQZiG0OYQoSP0tXSVDlJlx
RUNVJwhD99RcVcW43Ptl2W3XKBIXpqLcGpkUOGBXoOA7HDyBf3bZ1SnzAnnXLZOs/VH+L59/s029
MR8YEJ6yFUF0fvuiJ6mK0IvqGAajqBwtQrNZ3urXyvr3ImyP7c+X541j4awepjnCpDvtW0Rv+6yO
0H/Zhq428F2TQh9/n9pcxW0aX1jsKONjlsIZOLvhNl23sNQ2crKGqvjjsDKCE5QNK9FpE6R7BqAa
u4YZk+/U24NKMF58fNJgUJJDJM+Kd1594DXYbsIaFS3T5kTWGDwzPWkeYg5y289vWfxJOYGjG64R
UEf3FVbC6f8czEk82JhcA9GJ2pmaZroQI3mrpfK5EFRccq0E+W6k2rBcz364Tu4ChZENGIsDxOs4
rRqEIo7wwI3lSn9z5st+VbokK1TF3mQONGh4F5ZT1DxEDNKfcjd9ZVzuVKYh6kkWXLljsA+BJvjW
AbeT1MBNylWw+RwgeAmkELdQn7XflRJDgAuD/ZpUsNwQpwdyoqTVdneWtsVAhQPqJPC4iIkrDwW0
M/Gzz5Swe6uhKUDmH6unxPeF5e6gSuvoAK/gktDnnVxQuzIQIKL6q3cA8OC9gx3MMxII2L0VgvFY
Iu7GSjQ/tWos367mH7nMoCqnLOvpleE4kiOZ0f8BfooLYAjvGSbsGO8mL8QXJd+m/ifQhgFBo00t
b6RPcByRsB2eluJW3Tb2Zi2R1WHzpJT/U91jzTiGwyt35uyG3RjzoxyL0yREMy5mZv4oZ1U5r38V
dcbwExy0jEIQm3gtzsyhqXcFRSpA8RqMs6yl2x6uBO0/bq2P7fBXuOTQckDEyaQbNj1HwaW30f+2
hmwv8Cx88/7eg8ywbFIDtjGq5NcAVmHE0HWymcv8s6M0t/s6ArxmKWEn89HPvan1XMMdAvfyAR8B
DsbLcdyybMV3B4vIZqcz7Fey1hvG2ipi3KLcrUGg3FhRkyQiFyxYCO9xyIcPM0312+MDPyWB/xB+
d8ouNbcAnXDWP4tYUeASRFyCJVJDnvZZimY7t/okkVpU8lF/ZlO3ommiXAlZW7+wYjkBhvi7q5il
o+PN1EdFS2yK/yRQCh3M21Tx6mN//j8/yDZs4J1yZzCH4MPDBoSu+iIRqsf/oMgLDYXe9o/TZFBz
XD9pJY5ddhJWg96GZm0sBnbGtgu7LXhzC6BmOUIl/M1C2J4crLuWQ+IXwo/1CDZFoNGM/vk1Z4oo
4GC08VorOwAkuxn1CgInFGTwtE91hHm8pqEpj9YlMMeisryCu+3FG3qxMwg4ewvLFrV2XVabkLQT
frRg7OFHJmbEDnNeyBlMjJEW0ZO86s8F2QZVJYaa28yNvLtrYVeCZpVwl/fAjtbmMpa3rq0oIV42
ctvbFEOhmayZYA+kRZ/c9P6FuxMHjZp4i6Nna7ZLkFaIxaJ5uGrpyCJydeZNdtHBWdEBJiYMkoe/
pmQOC0J6/1iW/Ae1Wcgw0AC9jljHXO/B+BxjLlSUd+u17EMvPwVz6DFGaU2+vo3ohnSxyFKFFpwD
/6JlrSCuJB+2di28PKzdwAADc308IqxFaO6rMuL7COPaXvxiEYZCFfa155utALogdI5Jqt7ntrv8
Si2lHqyiDbrOdsA6nZ7YWg7MenfcwFdcV9dnwW+GvvIwp3oFpRl/K5dtyCiD+8CXgrg9nuRWgkBA
uFrPgi+AAGqlbXMYDL1HBWcqEQgpxo+9bubdc13jSBn8xM2bUbGlnT2LvSrdX9QIgvTq1wPTziRH
pMtfTLpQKprh5Cnj/cCRJhWyC2LO0vfbMPo2PxO/4+8SO2H1peMasGjO1F5PPeLI0K7QbXnABe4D
6r/C+JPOuAWO3rzTHKrbrZZxNdKoLym0JYFdFIVnBvMr5q60TbulnaVuu6MYFReCGiweVWF9ij1M
44VBd+JoJN/CbUuT6nF3KnhL8j7nNuXZCRrYznbBETBVBuxvY5XnT/MQNHURAymnkh18MesTMCGU
innQw7AaBiHzKv3BeHLYF3ehyVAI2kEMCFBmXrdnteoAZctRURq/OYqoC/z9bsm13MhRE+OinxHe
AUw6W+RchVmdRKJnhIOxQ55yv1O3bJ8ue+zu3nhKLZtpSsbbXs3pwwXuf9dSRTpmkf7HCL5q3ayO
leXyDpztEGi7Kf2SMB17oWeFS1GlovOMBXbcSe0BC/f6krXwGBMJLT4Dt5QmyHp9kg4unKegG4aC
cymKaceqI4R3Y6BZG5udl1kkYZiz3YPflPiTN3N29P4dWqFRzRoWspsuauMjgsPRIuKM3fuht+F6
Ay4eHhX9T6thvDOVdXIUCSlFMSo4JSLy/neEJEXqr51ZBMm+c5BaOfp9lUz53vkHd2GPH8AivdHh
dwTCCRJdeYR+r5D39T0Du9F3YqbWFYb+Lh4DmJTh6LpvYl7smKQ2oc9DWNmXnzVPd8kJckMsNMnh
66ROm4xwceCq+Utyp5tOcjJHf5mPPMKAe9HjE1IpvCznTQkxhgI2afJj8858ytVJRrk8mT8sFjmy
wwCfOwQoqrNHtjIHWsHRiV4bCHPJ/toJPwcNMmVHeF+/Ypv2tlNt0rAHmbiluguSUF+pWN00C8kn
QgASD+6v3GngNqhdA07pduMiND8XGzHOS36mijue5mFqO+aEDamQTx9FT4PBg3SJx1xKLKhyr99X
myXdOR/pA6jI8sansQPVL82tZZVDj+ug2yzRogdQw5ovG6v3o4E+Qw5O/3g2ZqRG7faRLJUmsyN4
SYZma3J32QM/zqa7c3zKJ6RM1I0YqHZP+vNEF0KGchryAUsR7Gv0AqESARO7w8YhbrJECEcH1jOL
vd3Sjw/bk5r5I2L1SA2Q2f3UhAoNYfXmgAXvFKzYakcLJAd6XndxDAmbQG+BAeP3UsW8NsNTG7Bt
78PtJWO817C/axyyqYdY6/8jeTjt6/3yT3voIR7EAkRADQv1bmhYBVUrmr6Vcg8490grtf7vWHbs
WA2kGZZuEicvfsMTfEFSZtaq4SydN5tHGDYOWjufem2beKkQZM/x/S76vG1c2CC/No1fdJhF1qeR
rdcXvHKlJjsPgQIMaG1fLz1XTBx/CfdxBepjxLyjs79+8erwhTbGP83pazhW/iraXHVLaaWwshjl
H/sEsbgqjmXv/pMSQQrdsl9yIFdVczGsJklCnjLgHZ6TykaE7o4MI/BkZkQk0Mjz9cr/4s2/ECcN
9saL/0xXhQ5CpflVp6j65DpEKzTzZStyAX/LzWqdS3+OXT/aqEa67YWEV7hhI+5xRCikkuRnIBd0
unDKq7CVnqCU0J1cHZalufonpSvs4k+UUuVXgnJsvQi7w6ICpjw+sEc7pOjfLsGWIp6gTPJtx8qE
ieYtMImq1b9UHdJZRkt72Z3FtpatjtmSPvAv0KDPxvX+rSKkwxWUq/2XE5iaga/FCmmrEfAxGBiC
n/W3hPQpwN/Bvlgso3MZ0SRKJ0/SmmUI/7Di2lvv65/qDaJvU3w7ZC/bmqVkh88wnnf+i66orEbr
XDar0l42msWN5+K4fMlNk3YG1S/CVuS1emLwoZ0UxLGuyir/ofvvgXwYcFvF4WAb7N1Fxj7RceVc
/ltRiFH64SkG/L+JyTurg/BEVAnLVKLWf7AwnfktCnGnE6iEWXMRggATukvL8nCTcRRb9mPvcYSr
jYYdPAD+WRtXVpdXOubnBeu9vPLtPKgvbXzkSTOF/5vXbCrZ+pVEGTENUezLzeyYwsqV5N/6wHIU
dcYCH0TmtrToeK7UXy5myNAEe/6FQUadv464pYC/f/gj0PYIWU9wN4mzaD9s4UTPiveEMwJvDeds
b2PoqU85EHQ30jvMBy0l9mpDSQGLgMmIoXvVMurFcDctZZ/QYLwZHlMqMEx9wf/TyjSEDqhQMGQQ
uc069Z0zIbG48wHRlif+zjB8WfMVhCXEqFoXF4hNKSsp9QE/ut/8izl2OKU+FcZLKVX8j8W5Jpr0
XFN60Hu0ElneVPRzpMs9j+GOvJjqo8p8/Teghjdi2WbwWx0ln6Z1SxhqVqCBq8oAwRBFNzU4fHWk
H5Fc4FIQXIkze42sXpzvEXUkEJia3SkPmws9IsnEXl/vpnL7DR7ErB8cEyScu/3OM69YNMFPodSj
lzqFVRX9L/sygHyoUcJmZzcEbdYWXqruaTxUVMgzHjmK5lvrs6PPrg995b4F2v13PJv3D+d4f7Fd
Q+HbQcaw0EV7vdH+hREhSRaQiUfWT2ZdB8MxnbKwboltGFYdWwRexQXGX5hBCk0pz9RnEi7Awdpd
j+7EKH17oLNJyjMjeBE/raU5gUo+ElrfT0YMqanngUPEjg2I2pEe+6fhSi0DH2/qSPEAJK35IPWc
pZ5oeIgrgX9izIgw2a5I/G7aIcCPzchY13HhVL+wzyFqhe8P4a/Rq02KDIdhJr+WyhYRduehItEz
o19Lzzx+idWZ1rS0qCllzp5Dr2AnTJSosADFgWqFNFT7xlb/prH7tcEw8zbZ6RB3GBeACXe956ro
B3DgmEi5cXHmJxZjpJK8BjW/GA6YYRWI0iokvGC9c7e6jRGsfPaxkkOa/azNTPMvIjQ3p4jIoCSk
zJ3K2vJw4XAzh0pEpyVahhH1xw+hbeCkrhQ6deHJM4XqSlkMf5u/5NRYcvBi0pBwXltRghvvAtng
vfJ3sujWgIkLuJyNVeZ7V5ifzMJXBDCWH2rBL3wQXnhfmJIFkinlizqq1Gurvy7hHhRwyBt1WDdV
uKj9lc7x5vTJ+p0zNZ2wHKMBAcmo0gMUrunQokscax63rYy4mQS0ggrwcr+EYnmr59enk4YZofVW
G4DWqdTG/GL6owzaSwif/HPs5c5MWnnRU2E3WN1O2dvSbXt+u32E4Es4iT3wZ2ogVqvf3OaCies1
zxoFUcgKys4grtaYTZT4zGXk+FDX8JKBCHrbGMTD6S0DHKl67Jwm9NzexZSuXCNI1jlwFBNRMaBy
+fkr+3vQrj+cL6euwa3TRHDdxxxseg3PbVKof8VqAg/SZJEcMRDcU+8zuGcMUJKpQgKOlJGkHtEW
rCDhN5qbGaGYKDhkOQJd39lWzFh70G3eoJ3e67BGgnhwOeR9SH0KYxFMIM2t0RyRwtMj6xdEsjbH
5biSq4VBBzgNj9rg3xMzCMqm6/eWKyiuS/AqlTLBsX2NU/yvcBM+46jaQprHYqA+vXVxV7NnA9g2
uqWaKvh3FsAle9QGtpnQjiVjugzmaIFYN9xm0zeuTBZ0B6pFxBWgIQLZCvQgiPJ+L8rHpAh15VpB
zlOBqVOjs7oyXRL6rkFzE9x6tvFgP7EumF6Gmve5zGbxNP+6/fDSvdOlFvCHAE4AtIouzVA64eY9
ee6HixPhP1t5g2j7zYYTobZ49cAlIs1RV/8PCZPDKjRgmkuBxtQM2qSSyCYw0h7XJ7mAnNlUs1ec
BV0Mn4MgcHwg9MT4Ydw9X88FLronLv9yRAzyoT5ScDQHF0+rP41ODvORf2TWIhqjaGVaFotfV1is
ufzOUZr2E7yo2nDInt2aP0jAYXsKr5Y6pTz6wXzCB4i5CbPw3FeMtk51snhvgoRqWC/7JpHao0zk
ltKtvS1CUkaz0XhES7laoXIpxNL8heFjpUoiAZGLcpSWHoxl1oH9q42KtDCaMPHQjIA5+JqNiCTF
yFwx+v64N+OMdVIPpb3+hD6r++x+G+xl0gBfgbU+U1RuO37xEnFi+IyRaQKzj122swsfHRLsDotx
f0N7hWVWRMJGKRobdYBc9WINT3M2kU5PuKx5DHv/xPI1ml4iLEVtIUHc4r2NNjw53isbRpUwmkqR
g27nSyiWiIVWeb5wpadLG8iRiFD1dJtfS0odiFqcnrVuh5weku60+e8EqHSbzTu7K/ye4OLobuew
AxAecT2U02EtxYlL6okcXB+XazPFPzqx47FH1yoioXxpzG0XVBje3qf6hyUyo7oQ1dBStDuvHFV1
GDqbfFy1C0Mt6eiy48HV1kaCE//uR68toXgt8erSMpNAWC8heh1F86PEiWZiRz+ONaIn7V8R+kC6
eUcIvZPZ9jQg2npbIW3CA1Cg7OBwe+mJ4zNZLb7/QfXbz18ybOzNTK9whfPA2EcNBrGxB1RjP26o
mLd1tGOAJ0Sc15cMF78Uevz3lqBS+MmKPi6Q2hvRr8T22wILsnKH4+gnFdduxiWuuNfzQ+K5eMee
ky8R8Q/qt99AhK3NDIkY0GXQCEuYV3/3tfEv6XBuzR5yJ8hxG0h3AUYcGuclaDpXg4SijE0vmoWj
pCSqlQmeQ1Tl8vzSaHAERm2BfvC+J9Xm9vthgpifcttdHWCExHtRkPRbxp/Oio2Ns38UGZuqAiwe
tc6NE3K5Y2AC1tgFrAclcgTjVrj/aIZT9rzc1xQaR1ZRXQRqcr8J7GtJYkNs29ywaVpCCBG1yCcx
zIFgnYVrfkr6tTRkqH5DRjwRCpaUhAK95fx/Mtx5+n5jr7gBmUv6u0CCyen36sNfBSoTfBzKJpeQ
p+6JI+TGPlIbpq1cYGbcUOSWezS3iqHbJqdKqNlDpCc6eiGikKAO51xuYQmbEGekoL2jVOupY2Qo
TVK1qLX7C3gsTxuESA/e5BjW8DJDeiTx/vVx8vbxh5c+lqBKvqvPOhgMvZtGq0WoQj525nKEBR6J
1ARnpF/EIgMXcfyeK+DGjN8XNtOK2bue9iyaDl2vo38e4VwT42Uxe3BjSjPHmr6XMFJRmLbXijdR
85HPn3E6wZTXc0w30g4UezUUSuHryuTyHAPcH5JmJodK3LiTsvxOPztj1e/nsRagmpVn87ihihCA
TifNOVZX32Jwf9ZLD6rjOv0y7eBzzcIcisf3cjHB+SOGUzXB+UnILebKCgQQzLgxeGTp8M+ovLMj
OmYr+HEUaHmGna16AuoEPH3NI5MGoa5jmNjTTjmQuwTNnFTtLyfi1QTlxHA6tgz/2QBYWj5sHCXM
oM86c/0ejjIKdLFqAudd3bDtvV8+aYXx4zS/XO+OxOYCpekPzRTpwQc6dzMsjWHKb6jozDDBf9U5
7uL8RQUsQ9ghagG6GHYHOyeEaQigKFGuMZenAAlGtrJ+o/3C7GMh1titqVWsi9h017bsfawmi/Af
a0EtHv7/IZ0T3ilJ7+Fxi2dfmJ7hUQMdChM3n/KxEHhGsIxZvEVdNiJ5KYdsi9p8q9B34fnvBRYr
iWKOsIIfj4lkic3ZbNJ/7QlLUjReijbSM1lnJl4YEuxVJmGnzaoDfLkFXUfijPDYVww+EweQ7fUe
Dc2W1XEGLpp7sfzHd+Cm5+Ll4fMsZTBpLlMUysVQqOHW3JY0NJakY2aXDs02EKhvEqEmInjhWArS
WU3DkZ8XtJgt1wd3RS3HXxbd2OfTcoKFcN898Iglu/WofD2UlQ+NNgsGLdwBQJwEa4l0qOYFTsI7
wpspFYT/VYTYKeXeEFYW+XHLHbr1OdaUK6MkSBBC6At61XiVwdj3FSuLgVVgR2N6h1MXBKKHSCvC
eJNEF0wnKXkd40f6btZQBKEHWa3ZklTaINOqCWQ4s73MSYjTHxzdmCODOvzR6VXtI1kzwVidZnO5
e7P9uFGQkSd1tWBKeGbxijs07jI0zd0rPnMBDDgQuy414nYp/kVbx4N6fRXaAHpO6I+ukDUYLfoB
5dg06G8d8lieN83HbSB8t7YY6IQcaVx2HwdknZvOzv2+YoZqrNNsMZLDgRzw97x4LwVT+jOKXnLZ
bYR2G6wB6JpPmGlCXFR97W6Q5jfecPVTq2eyZpE0Tx6ukWPmaGYESJeiBUjmmYzhJC1ptKgfCeOW
ggScvRyPJbJZ0XOLk9ekmpb69vGCVQoOILbJrAwK3eodsCTE03VWVZyzHKJfhOsCpdZ/z3VBz2hg
AvYTAkvFdWITOOqUqSzrdNxQYmOjSsEThce4p54VizM1cVtXES91fXCo9q2e+AlTo88TRGKWQIPZ
DATf5ww4RgwwDW/sGzcdcVt7PQHg6j1Iiz+OTSdNov5rOjAiyr69sLDcUToHGGN3L9WWEOxXbxRY
hD7PIuS6eT99HB4g960X915WWNAfqWsHfzcSyYxvAprkubRB5b2uuDmd+D3WJbe331EwRYxvwtCy
pylI0DL698cNCIrscpEhSJi+dv9ACYcp3YBnlwD7yl0YI8KxwsjzhWMsE7YinyUBr77kfUqKi225
G8ArjjSM6479bIbJA8qfKu95DWNAXtnI/oZ9An7y6ZeC/3r02QWES/ojVD0b6+OtWgkcLkbiPK5w
X6rnf9Q9eOmpvZXc6wEp+pGsUl98EwyA54jRVEZhReppNkUMO10f6dqnSp2XdH8wXvNYD+VFYgky
RxOfybvpVhu0aphceahnBm97hj+VzfFxh0JpyAKtjOYRvDQsMoaewwtANyL66CPuEUTPY5mt49Z1
bC/rAdqaXByVgpWrPawD35pt41LsE8mmC9Jhbh8Kl0A+vVLlLnidGv0PGzGE0Z1+0PdjSKOjbEED
a2G1BP9hVMUET3IrzemP/3k/JSQnxklNcBEROn8TTVwOQk04FUiiaIQ3nCyCV8O/4jZ7qIVXtYbO
1LgYQ21cLxRZNgtpcpteNfRZw1DaATFHZYEPXqYETOEFUqJV8jEQ0fawA8Mqu5HbC8HMDYXCgShv
GYEKN0t+6O4dWgUJ6zJXVI/gg/eU0mOUAWSEQ14FY2UIlMkw/njvghfQzJhQA1EoK4YCvKeVToqr
THHZjoeQ3rscljW/rTZJKRSY8QYbQIJmmLwGIr5YghJN0d10Xob8IPb7hVNhfPagSj487vQxSsoz
1AvGgf0YapSMrnOmXbUumRqCNFqQlXKl3cBXEpcqVjzqaSFykTTYj6ZVhQJvibEgIdnwWontJKQ/
4PZ1Q1JbvsnbEdcgHvuek1xO97JNPzFNkkVQv5qX6Zwq+5GrVYqpM5KoL05e7kgeQ0EoS4FWvoDD
51qZLPhS9RvaUe4DX2i87krKR7qK2DilrbV+ccliZDCmqXihC+Z7hVMn3pLpo5k0c+EQo86+6rYG
3bnRQaM5wmkCtMB5FENLfg3Y5feidzevHYd0iqWpP/tg+yEerXBhokbsfcvhRdEMqOYLskuSIkV2
NI/x4Jn77sQX4Sy8g7kXlVqoIsQ5cJHhvSnnKV8RxummRVwh+Ztysl8U3cdUkkLDcdAmV3bO/iTQ
IcdkYBCnm72Jm7nHTP7u1ZnwhmUsMaVshkPKJqiAtwYBZ0G2dpZEGW6cv+lQEThlBHGAOCPPtviK
9IerCFGCGiktn+9Q1UF6iNwXifEzGLJF2/qW0YqXBgMD8/r0I9BezYNgxEAkKib6DX1uJY9oIEmx
SN3Kmi3B4lj4vMCNVpCMTd1ERD6pVFW3TjqlByZgCaj6bWXH+PtlXGsc2ZJr5YTBNwwQ3aWwVjZv
+knCj02IShKK6pgUBXrnkbsNnn6f8T5YG1pQDUdHAuXuN+yn5EmFA62+dXPU6sZazJcvZVDwBlFp
VsB+Gy8hrX2anVa2x5F4UXzmqeIUWBgkqEUn8oy3zj0O7rGTM3GyeJlV7Yy+C60x0PQmI6i84vWC
fZ3MmlnfQKwhFQI+K2gciKQnWyCYT1QuzkpZ89DNfmckIYDU5P1NiQ6PwNbEzSrwTY7eWkAWRMZW
oCl5QKFgRF1oad2s1i1lSgj+0CvXVyZL3H+2NuGdXPL24eehZDtjil3VOm3HrMs7qyYKSg76pBbm
kPsqnWLQOw/Jquoj1ETR49DT37CtiQ9Nxn4PFTdeWWkun8t4Ul4xn6/2Wb0Q4sckhNdKWuW8dpC4
/Hx6MIQaFAhjQ4KzpimgU6r9K/DBRYzBQ4xtytcWy1Qca4Un7reDciRltJKeCYDGAqpGySq/XFaA
7P9pkTCYQ6IvVraRMWLcicLNjQ9QMd7D5adyYrcLam4kTnNSPCGEpuzKyyvc1wRzUBQoeAhe+R8L
oIfQwL66qSB5J8Zgu+BSfDd9tuxfgFmomtGRe/l+aiBg0rpV9OGmQ3M6Kz08kIpSUhrE8DQ8J9IS
+OyiYfBaG+AQPyQFQyzD0bowvdJ9IkRmOTFyLE4+xD973/1Oqff2EGt9tW3JK4VLlr3x8VE5JrM4
YKmRvZ4CWCCHMqjqb+o0K5rPsKfdIVH7Ep4gNou1SkhOSwZUKbrxac1GTLDtWxJUqVws7M/ztEII
H+55kv/9LZJVFbgL9EEIhYN2xSbRh0obB37k3NbOIKO182lPNvJfpZEuRRDg3T4liyYumsmy876d
pBXXlwHWVR0Y6dG+1GtPL2UcvKDb0nynA9OYrvNSK2AwV6h4OqdDL8+vJLvw4/mKSiBmi1rDfoFq
B4304GTxgjphNDGQLbiYTXnQxkqLOD08kfIzs46xDRfOBXuMjFvKzE6nCaDSNRHb3CWBbgiLgqPk
PPN2f2GvroL1rr8OC+0mh7A1k7GmVxDtx4tS0JKRdR+pQ7T6+qGQ72ZHnryQFd29Qsk5GtYOyvAN
SUSAHJt1PzqE6aKRlthLDFUwqHLSQEsos7mvTb1aRnzmEjswvKxEQaQQ6wotjMl5o+28brOj2fUt
iD0l1TnN+RMD36o8IgWHoisqU4WcWieoV9qzm3lfe4pPO6JtpZnhQ7CqQG6jo3UdNz1E5VCkkWBG
uU61W1Jsz0h0zWldTDEUtsxa9IFIfR3kD4kC0i1LvpQpcxsvIj6fWeNqN+RWXxmxqvzLoVkVH9CH
qp2zYcQVGxZSzXNW6CTyBukd6l4SPz1E/EKV/HxPv8kNF4Kt4X37fcJKEqbBsfIc8jMY9AROVXqH
R0pqLvdkbjqZjs77zc9ydhF0JmgIFnbVk3h79XxbXuCs9eJ9rpiFfkGdYVLFRVxXa+eOfQhjQpZ5
5iUEPkTLRNFvLZ3pbkGnAjCFe/+qCpqMYpqYK9YcF4ehjIcahcXMJlDQL8erx0krJnHl/pdiijVm
QtFuQafnIQAeDQpyXgsISqUN6vCelOOHsWIs02nAZ24HkOWpfeBXuL4MnJAa0qQbeUX9FCKi+ovV
F1/vulRfxX3asxmah2OHsDqf4Vu6PrKLplT5B6Gss13MKXRePX3+k9I+3HnANB9fIsUeRR+iOhML
8ChquVUr1c6wXqEmde9Rs+ghjxW6qShE8pc5czVKbHeLO+V+1L/AJVK9/61qDg3rJ8mXsZWuUMH/
yoVayAiYJXwBCuvdE/2qOgOACFiNoyWTPk6KfeaKEvz4gVYRSJNYR4JQDeptoUNI/wd6crZz1UkE
AoB8Af+YOfxFUuFyyk5wCmOlw1qMscIDpvhYVqC0VBDrU/uDdaGs0+DgH5im+aoO5iQdkOZRHuqe
tdv+QBDAqwZd7QLPJKLYtyMLeIHE3xfgjU3qJr9MMJ8UeCGWQQnZgsBVPZuIQ5jailYMkiL7WXdb
HUbkqmeABX/f2MfV10lKQ5xFM3kOr9juD0yVtgPPbWP7lTXKIWMyu/DWVMpp+M1H0SGYDR7mfwRf
PoIfjip2UU0DamggC8nv1dsa1dm46IUdSKmOz5KfEiitNWKh4NU7OCaMKtp9Hdfzy6ntEBDD2CJL
/ACPp0NLY6r0C+g8CCa3qQWBf8L8tD+ZhUJdKQNtiWja76vJfPPMED+DoDOv7aSbHGbCylIEQXRS
fQW4s0Ux55l6XliNuVNcQLXNo2mfeTM6/nnMrdK4k4paTjx9LrQb2UFQzEbLJO5H6k3Cj0e9lhiu
HYjB1cEl/CuRexlxh/9D7ugh/QmwfHxkyU9Mq9tokMpk5pt6FINRcQTR4JsMUWVV9vfdaLLjUqSv
hf4bVSD6hkePHGXu69S778QPXNii22Uy7QWly+trMyQpf/JYkTdFdEPHSrd3lcYOZctA8BCQR445
73oWzCRcCVHFDoFXIxk9XhjfVxAlXRMJ4vB1Chapfvdrr6uWYsHaWQzziNeYTC+X5BJqq758hKIX
DvMnQZKgMSdeMEoM1KnQePn8l3wJ/yg/JQJEpfS7BFmFPD9P8HJufVr+1866KaRdxro/IJHHqjG3
yWgX7gaT6M/4yoloWUZ+K34c8CFjc8bYsdFjVI01dBGtD5azKxueYynqYjopEeK+cDb9ooNqY9T4
lcpQtSmjhOAaG7v1rF8up2NMIGqGmMEXpbBFpRtm0rpLFXxJ1UFx1Ou8xj3vl6SvxfPtbAMjYAVU
f46X1r6VC+ulu/x1BcFYkTXtRx4ytvpzTxbHuMfY6mnq7qjhMAGk6yZgg2pBGFKIPBCtSNKh/oII
R0cqbSLMFWL6z10WaSSntPihW4db9XcP0zrmAi9yzXkJDaU6C125SGnXSVwoKOkUR9fj96ffwsep
ffrkeI3xsEnQkR2bz5I7KvwptFustRy8mlYyCkyEEDH16LbT/mTbdOoeKrPEJMqmPkFKBNJW/zyi
ALcMmP5XK2LKD5oGcnQwKMP4PwoXxtSscYZT7t9sohGVpx0aYn3moxXb1xxsLqWdO/sJd6lPFXtb
iuWEKAijlfTQdCy5YrtMza22ULDcOHEOtVt8c1psTvo2JQnxr/zLOSOBXnvdVgh+EL+acnOAzMfm
wL0ht7JhwYmSwIVXT42xrx9mTsXokmNsIxemeVhrGS5TV8zE7hkp1gfjYEIgo89R8DsZk7zFKLUJ
AJfOqBbWUBJ9ge3BjZS/XnpEoQMqfo/OhiuJW43HuJEB+ixUUQsuVUpH1VU1/u29JZVYoU7zhqqk
x8QjX15hAnjugIS+d0JzbnCTX/xfcHxmlpL6G0tT4GN7G5KJyVY8gxVl+e24XiDZagHMhsQNSmzR
YVtHPr0C8LR1WB9vqsMJhvUZuxukqWbfadA+ofO0ow7jyT2rP0O9EL8Qfs7pl37sSThzTvtLg+Kd
lPZMDngFQaCbrdLQeoD0lHlt9GZ2w7oQ9bY1Lx6/V1nNyMXGnzddwsLcZug8jFpU01oXNKQQc0g9
AUFh2KeLUZqwi7f6oRq9rMY7GbiOcOdV1OpWeppMHaQJVuhlzJjSOQ/9dDN1fF7Tvi7rt2nJa5pz
e6iUp7Yret6wUcHt8h7EG6uobEmWWYIF7/R1mald0PLurul3AiF9v8TCSpfzP996NIK/Vd3IdUVo
Ap4NaAzWvvNuojdCQwQTlmah7Fe6BAufDkSBc3fSim9oi2Lxl2WM6uHBGfTTI8Jc/4+eYelgZXti
iti/DFMg5+gq2IyYUvCUfSV02MC6KWCXvB+MDj0jZNEo5QUDFLyV4kNEWrCEXEBegbsJmuPHdQc/
mMyBgqwVjAowLp0x4MX3YO/WQySPXopd5+VaBMuv/yT7wIpPzt64vWDzOHl7xPNx7N8YdLNkHpbL
A7LLLdSaQnRCFzkbMTYW6OXDlYKIFiMRQqEESzfM9LdPr9D+6pJMy/5c5hODkQy4s92FR6j2u2fY
uUTWbQ2UH5/igrE3TJHKupfBsoriy5qM7NijNycDbkTQJGArzz4FBvshN08JQeamtekmqaPm0Pbd
hV1M4bG28y6hf37N+CGgU8bFfBhVrghlcb5aVcw/8BZa7+A2dqYa6iWQ7PVYdSVndINFLkfnuaZt
XEPGtqYw8QrkDZcF4qJ3Qkp96KMtKTEuFeUB97Dd10rFmoniDeHhAxA7BR9J7p9kRvaKyh1J7L9M
D0SR44ZqIhkww5pZ0TbG2thaqCyZfvZpE0ytcl9cdximdTIoVwcJOYS4LGuRO5JyfSdByDg4nQof
0SrlhvHNYojWrGLuJanVHr2CcSREd5Cx+plc/gFcDjA6urjguXX+7rW4dBQjZfoA7CUqldz45I+w
4YY1nMX4wxXeIpoJVegmBV33nxIQDWLnzWD1c6VCSNjCDfapLhC5OLxe9i1Wc5bJbIFub2M6mKdp
uJ37hB/Y1svdv1//UvZ2i/by7gbR32k1FyEf5CSyJQ4gs/Z8KHDGLee3AQLbavvwQs5I4HEhc8rq
l4JC10QilUMdyisnLnd9XgDbxJySId+BGIyb1DqFXGu+7DTicwevFl4ri49/xB8dvkbKbr2qcMc7
tV7VncHCrPA1hFdoUophdOya3lHEvCixQ0GgPpVUfBk51qKJGtt+GYwD+JCtaxX8RSBwrs2QOOz3
M2RX2NmTS+HyOiOGP+MKQl+YFHtp726oVdEjkFeK68XxG51DBf1RF2lEpoddnBJe7e4K590cSUZN
vOOJ6on8pdQpoODM9n0vfdjC5jGripcpjrjwwOjwW2CqvzmTHZVweEekrWVUTg0CLQFGw9++Twy8
ES/8Egt6CHmUpneO8ZFpkTK9D3NU4UBK01XHw1Ml7/gt/FI/CnwNgxRizYXrYlrFgppGb9DIzCxV
tfehfQVBumGwl6sEJfY1rYGI166fv45KBrXwgUXNZbV+Dk419ggpJRN+rblTkqEiHQkjH0exzVNm
J/7MR3KWBCTXJQNG+9Z2HycO7jzpxZjjw+8EzZPldnqMZFZ6OqLTpiQQUspCVsjRpinrbYGT9QQk
qjlx4Iel75QcV3r2ZHlmBIntIOZ4aZ3hxIqlT3tSP7YsfOuFV/xNcMjX1rafQjPnSVCa8WxHkAKl
ysuaA1OFIVbYMzHztWEk1SJNZZXWmPisQxSJ4WC9l30I8TZ8U5UridJg2tEWxSVbrg2V0wvsPmJt
5+mTOJj6T1yc2UB082ldBPE84emePFL3ErV8iACBKvBjVzHo+mxNE5+mP/czCJ4tQox0Vo0jtAe3
82CbNg7J9Dpd54LvGjUZM7PUFoTARlXFbnPB4JNGwtJzgYoePRklvunKz6nWSU/scjLwZ0C4oAY3
93lMZRbjo6TsnYjDDf6+8XwqD5o2f0aFpfzqKhH3i2FPfJpUxgAWMJNAoYY7mo2uacYGjelRIESL
ptcJAvAsPJ4yepF7S+JG682a6NijkJqf8CfePEsFucgXozOnbkRGFkuUpD3iUSUacF4ENqMONhho
v91CcVszZwN0/4ETlrmPHQkwHQ3bJm9BejQ9uEpRfBfGj1Zr8RCbOqNK8PDG/GcXirJKFEL7UcVi
PC7Ae9ohZnXKsqbEkTsCf0NFkH8hIOvotroauID2dwfPTB7ktrvFgQJP9bwMadXwX4HCGEt6+ni0
MU09uVnPx9ro4vfmsjkx0ipmLUPRE4CiO+s1KLGTbvacOr01LxKF6TXlUtz1T7pjDBIYDxUUxN6Q
3crU+uPHJ7E+YIUaJCtIkPWjYIu21a6tO9+J/DJTK7cHi4Rw5lgQNc6xYbKTyR3mFBJeUmDJaESY
z1g6iaUIBz789RQQYFPGqbms3gDmV56t4FweH18D8/7SEkgJgSs97pa0bg8z4rO53X34won3h7oe
81h4SYNEWdx96FiaUGKpGXEOdaOVf1q1juAsgZDpeXXXxc8A8AuL9JwWyWTlGNskp+YaBoj9MJgZ
UF81TSCdgVB0R0VCCD7+yjIGz/O9Yf2W9T4BBD1ryCCaB9kV8f8KWI3loZo6yVbReS72svwL8R4L
ex0kXpzhaX5LGrZVSDgXbFktwHslWHOi6K+DQ8h4jxoO99B960AairsOr4rjlc1upAzvsaObKM2M
huuCtD/9HAHnX+Yj9YE8FfdzX+6STIuJuhrHlhmVwMtTQS7l/yQt9QeR1586pQ0CHufqgHuXkS/g
wFGifd9ejjXwnnLfRNbA78JeqLW2mgxEHsiXb04f6idfkl9NuSBnVinKHB+5DbypD5dcZePYeX0q
6txEAyGDQlpf41ntlOrFPrQRrzpxWdHR6Lc3fh32U90+99GTD+mttwmcWv7cVO04THdc8jxNsc7s
lOIrPFBvRk9BTXsodAguBI5ONxrE4WjuqKj5hox28EJSSXkJHx3fK33GqvYLWhOBnX3HIEEEyBlz
4RgJnUlYbKmWXuC8Oc0x4nAfoGazkFMtR/6NBFQh530PuP+EYfLad8Ie1c9m/muRbUFgcdghkJsr
fUFA8YqGH4K/e8OR7a6ckmLaHB1E79K6LLHtg4u94FSS66h2XvQhi3ICmbdHjelJIUQX/Fauvxrq
mVpOxQoYQqydnz6XZHeOGgzq8IAYQonqOGQNnXuZD3GB/Tbb8yzg+8F/fgEJ9u7yuMsqL/g0Yrvk
6BYhSu0r692J1FGDMyqIGRIrePnsvynoB8CmZC9mM0FLbHj/0hYPrn1qJtg7levCNSV7zVWbxMO8
SZJNcPxJ1RbEIXymUEQtlAX+265K2d3kX4sQB2iyN/HaA8sV9F7kez9T4jIzJC3EqIY8+Y4rEvci
jSWvGiEH4In+2gElWxH5NJNnX+Nhk0F0foLumhCeWIQnn0hu60qW0o7FiLdfDrb36IszydCtbAaL
8+dsQrcJvjG+39/xFLcFXhbsUWWXh2lUodwxlZI/vjlCHfWEFmy41iDIfmQmDegQr655JhozW4CT
WYpedRdXnTUxyg5Xgi5K9Q7DUYvOVpE+5JGrsbFbmK5cgMA/3uTAshViqfDtWFbIniLzlQeCIwod
J7hqhLK8pK2MkvPyff3NykLBfruUpxkMiYrpY3t7uVCIM6EUIh8BcoxjJ7ni9C+uc7ju5Gprv+t4
iW2vVqWjzHvtZI0gDLITlqMAqpd8DvuioB9rLiES5i6LjhScTmo/7KAsjDOc4GFgZeJ2sMJBe/V7
H+X9kY9zAxLDKEVmDulKXk3Mnp+OL8frnD0ig/EVQ9uQku6N0kZaYgJKvxMaoIALt3tWR+n1w5z7
jVRY73cyUBCoLw0fZCkw8216+Go1uSBHIK54v/07KPT1SGZUjnGihUQeZnjhGhTVNsb5MOVY7wPm
0L/jd001EA7NCyo9eIJOWX5yc4u+Clw3lfseOjR5VUt7ws60LS6WmoPNJEDZpS9RVc5g5IVOniHG
eCz94nEDCp40H8qTDRsu63PPFEQOw7PCDnnJpG4wvut6uIJs78+697HEuoLaJE59E7sv5+BOZdfF
4Bys6631nKcmmM7lKsta4mezzG5cTZCE+Jm5/Pyco4P44+Z2+YKc0H4wvmE7pgOCO0fbYVU5ILW8
5mWkoaElP0QJZhh7wpb0LCFUuqtSztwPXEii1btaAi+NbHnssg4ncPKx7zHqbIO6I43um1Fp+CG9
K6OjuA72ieeyh22Dh4zJn0hmKkNJmkF7Sp6g650cNvGdKcdSZWM3C3l/CTtLMXPYFathZsBPia2A
3DqHP4E2aLve/vF0IIwHte52LdY2J93E4zT6sBnu2QszDLAH+XX/X7HygQwR3LudH0xdM9wxS9yf
U3vcdYf/589dW7p2/7UseTZp8GHKaP31uyzAbxMBJfgFRUQFIz3ktWbRCY2WHc6oiMJJ/iND4QNo
zS3Y4ikRq9tUrGMUxz1KI+Rw0FTjGmBGAgitNLvm/3Pl9oPpJY47D5UhWIbdahjFj7s9EeHyWIOn
Q1+/QCRHwf3R3pU5PYNgv4BxgB/7JrbSfRXFOePBb6+47BfAjNmL6m96imotKdF5mpSBFKZ0LR0G
ZHk7/8PSKwokhj9eUmnaSddOX1oTg8xCesPz/I2s6pYz2UQemSxJIk1NpZahvuy9oRRS9oDSc7k1
H57X6M6w7Q0NNdI0tqiMe42/7iFSwek4BAw/LeTqCDHa1U+EtPmNTyxhvPOFrfMWNtI/qIMZS9fW
H236OGDzAqsFQk3Qfqpo5qyuUZB0URBU+udiHME+IXttX4zuhQKrNFjEjJ3xpqc53W0rQvTY0Lh5
/mx2jpYY7LgFusyOFYIOoo9SKip1Tt0elXJlm0WWd9/2UZI1Cu0rYNPXRuE5yigsoz+XFCdfjbZA
Jh4DB6bOoeQxEPTlqa3RtzCIb+yMVu6ZtQx2StoYN2q7ogMscPjIE5X+M0h4EKOGe0Yy9QCJo/Wh
8JMdB+EyQUg5EQrkb1BA6Fux0oqLO2E8Z+j0xOlYUkZ9qdJs2YhA7wb/keicZsPxspkxzpZTMC9x
opi5tBYoRCOZvR7ztn4eZ265d3xqqWBVMgqCOe80g2E/MTXcv1EFVU7PzIq0eTyStf3WdJjTv42U
SjUBqfC+Btr0VqM4w0yrUQEcoyEl/G61oAA1uk0ADmjBsKb/k4m+Odf2z5dtNRSPsMswf7puFpXB
zRTb9saOF/KXX/5R1ZvK0nAZVsskhypo98x53nQyKrDmVhxvftYLn0IKbL1/iCNUXrEE/qDgB+iE
+XOUHdALvLVum0V4bPT8vaMTLLuumCGTpKmWiybrtQElIFFZO0K4mGKih+oBLVt4JAK4CgSRaaKV
4Jp0cC7Lw05A+DUANPwJA1M+o8WQN1rEYjnv6xJt13uT05WjGn1DNIuVjVsiRkSHLu7X/JMJK+UT
tnEpEvnXNmct/RBH/+C4QFQDTqomPUn69/xOBtj5LjNcGx3Cof7rR6Xs+SsgiUXKpr+0F1T5dG2N
7t3J5qXXX/vMwsBo6pdeUsAzOo9Ce/FW73XeuRxYRP/Dov93Gw942i5OuUknuI/hpGV53F89cS2l
riEBTeSvS3/bWDK8IB/KJ0d3j0EHxIbIXZEVzmz83rHxhMEJj5TwuCps4kr9t7NI3KPEsDPDQrmT
Lcms31jTCpeLg6CB0jcCC/zGHvreCGXrO9NB0pPC3NU3ASrw6lGtBL3nKNPDynk6kAovw6en3/JC
ZGL1QnliLjonh8+4I6ndsXqldNXpCFaYE/gCdv2+ypXA5UpVTho/wsvkDbOnzKOoummyVDxkehdW
8czAyg35UWyQi82P08uuMAXuFtwmjjLm8aX9GgGvXA9eXqtAO5UGI0Ds1Ied7Jvn6BHaseChxLRz
dqcudauKbmlSn5vSBU+sDz8qYyuY0lHAMilG/q9a5o3NewOWT5MMHrW4UC9Y1YJ8yGo1F7XQ4/K7
gNf43SG0FXJm1hahG0nAyv+BmJVpsSUlQx6YQ+CsEZDYMtPdoYDClQ0sbEEfpWvB1XNssawBcsun
yv/eh0uotPIzcinz6LTrqzcDCYfxz1nncMvcdM2XEdO62HtNWwuh6q65pg6VL2ClwvdGuDe2waOG
2tAdSfFZLOotsRRIhVuFdBOBRXQWBN5HuhBEH4omIEfBdBx9dQ6ZeYBFRdLH1k5SWBqA3gd1t7ms
zNntxgUs1UeS0PnWSLKnrxt1/Ypagzv/8FbOS6ldYHtYfH1qKgN4i8wcrW+RuXpPmHz71v2BXGUX
NONdkBjGiLhcUOtllJa8k8witoA9OddKpMbYJbOWkK4fX3jguAT9ub8dZWAZxQya+MfSEEFgtGln
HVQc2dmQN5+hRuku2QSZEbvES8aXR23Cg9wNGqGqZfJ/hmC9x3T2z8P7H3bYDyoiw2ZBAQH922fz
1TXHgkZyKgj5PIZhLPlauOuGaoirUHmSkNhN8faINPUwze4mK75jpkECIkfiDiQCOKARkia5mKnz
f9XB9VtU6rVgr6XqcXc9lN1qfSzs+UQYfumLWYtG9yy5XGBPgvCtiHTWcxcBgYgF+7qo2BCKMbm3
D9RigG5Nj6uoMADf9WkoX6rTT4N3s+P4/JnHGOGxJSyGV/5StHDc7urE25HW4v6W7I+cHKbtHkGA
1R3imbmVfUBICYuEsXftTrIDJODzaxKWG07KmeBvAWTwo3prFcnbro9b/QMHZCQVeL6OXMgjX9WP
ZdyqiCoyIlYkyu6Uq+9+hESmaefEOCWPSy938Od+Y95+U8C/SSy334fQKvSesj1BJ4KG8KOtH0LA
hZFuoSYY3XHfkOP9e3UVUUu7ibWlzFhi/bOIuMG7i+rKSgjxDBtEK9K4LE4KuEHAndwkGeJi6pRK
/iabvPzfGKAbbH7gE7VCIueQ9upg8zGk6ZXhXEwmZM/Ic0JO7Z4QO/crBCVl0+6KwywGB5QyXCcf
C7UpQ53ozn4vnvqgW9G1z3sOvezOPcnZ3BnEsMQ2neaj+3O1a0Wf2fH7eu+iczyxVF+MYFxIUh/m
1M83nFhZg7aMHAUvkYtQABjPbCjm7A5DDQ6H+sEMGSm1PLst5GgrbIwOk2lvETvHI5nCX9ESafm8
+bq2B6g5aTV7WurqCYkVXl8NHHRMidVlQpUqRHLpIInFhOuvVqCL82+XsvaW34Ng4B5OJPLkDn0R
e7QXySwBMsHY7VSa90zxzZt7AnggQ5si0x289MdnGtl2iQ3aD1HXXMd9chP5KaVGg3Y49Nsf/Tpb
27iyTaiZFmej5y7AFqO+g/SVY2kKQzWDqqL2QNDMd7aLFL5DmHEkoQ63OQyzOGbdZWMQER2KyrLa
GHADCwCylttKD6cSXM3iYntiGlZZt9IrGKvn2xAEigcHrXktbrF/Fwe/LKmbZX3zjzufUuwYxC/P
RTnEbTzL3eNAUzRvNm8CnYU+vM9Bs+ex/258rYN+CqJDzooGNT57OmOwKFddw0BaTyD8KeStYyno
/Rxa3CK+U6u2ZbxA8/++Avo7TTMm5Jh/X/DbzIZnzh4rIostIPfC9mzFY/r6Da+PHQtlyC7oCTVK
nz7Z4WmEXEZuigmeS3uDlkhhRvOiKSIjhREWPAckjczxwv/u3j/eP+MMtAAl5ndnwj0o4ARYmBKM
S7mL3b9+hm1UglSqCjx/ZYR5k8a94Gy+xr7AhTFFQFqpw/ZNJ1N35TiHPyn82HkAWK5sSjWEysEv
7XkVeMHeD7ppzgzp9upTCAJaNWN1QGmdPDVlTtV91cF1h0sMeoKfHQRCgEYrjXfYx9SJML9CW8N1
HrNEtwepZyg0r9AJ2w/N6HilR8akdn8MZ9/yn3tfHBD27n0rUNUENTP/A8h48Jnze+2qordU+i4F
o2zgkdT1dBA1Gs2oiXLHgLpzSfRAtiNPDYfT63kqOt3sO+ELeMsTrz/sY1IghSfHOOHfy3kQmbSy
yGWDx1QwrIO2MvFw0tvK5fD6FhyuBvW9Hm6hH38F0X0iVzkW21JPGdXuY1SQmffesu83pw/fCjds
APDWQaqDQd9KfdE9ki9dbNH+js24EnI+cEsN+nOjqf3kK4jQlb/QZThKJ7ZkvXUr05TDStvju2I9
dabfiVhljStdSdPq5TG4S2yrUnkTVG7nLYOZt1/WqrCNA4u1Yqk0OsHRfYrdh8ikr2J1MaBl8v8R
mGAQUkqtWw6C8h2WhOice7qwwPCtFufxtjMZXktmjn5cSAzQulVfL2DP+xJnC64M7EkumtqwoD8u
PqxTuxmH7gzqVpCA1KpwGeNT/Zd16bN6uFOYgofgPEDhkKzfVWMtdEhLBpkuEkuOGUvJSdLmmLTl
U/72PTSbrRFiecRKGuprfqbb58kQvnMQnq5MXbuinY5uQ3Q3Ib0D32tP9kAb65MOA9H2bjqMqflv
7xaEzOLlPILbzYdB9FhIAZummxWGTo1Y2NlEMfNwG2rL/Xtr68a/VANXrVAAAsayHQcZSc9il5j6
vIcysSmHPm3vFqYsiEpaAm97wvGOgvGONoBUR+SP5NmuJ4CnCSS9BnMQAkOpJRCPfJMAvebcPgJ5
XQZu65FTnwUHofCM6hRqmTB88oFwFMVKArmvRbgcVb3pY9jXYFSlIMf6cmJPebGBq+DyWKRkceMs
cb1HUrt18Jpf4r5h7cwqbe/EQpTnPKjjSR54PGQZPtT6HX/yRJGslb+R9ddScbhDVpKps9o7uRYR
C8MelLeg8W5ywcQjNBURQuL3SOpdUPXpmchI01ZlpFV8uMBJlCQf7eMQ1M5CYAg4lHzGTndrMAvZ
rUq2enBr5gBAtkCUvS9V7sxu682iJ/SBrJpLD3Zo6hYTvfBzOIP2606UG3634OouB4C7F+i56ndk
/jHmZdVUG5jyTikO99ImMjthLJqjZAKYyG/mm8CxRc6XGNpXCP4eJu4YSLNmyeuTxdcjVYdOEIjF
uuVLv4F1NpL/JNYrfrQHiG8CHINw39gH+gxZyNefbqB/IpjGbxyog8Y1SjwqKU0pUB+nAIdOMvaH
go8UaRkZKhuU6FYHK7KsHMJiujOCj7XEqwaFWjFCO4wCGpfBWb7P4ZNj1JPF+w+WztFqdOPi1et8
pR0TmjsDn4ZRquhAy0VesToLFLNBCE4NMtxmM7EcShlbU+5xitZmEIump0OQ2zkwr7ShsRPgqmnu
B1SZ65ZEufBcIuOi8/aP9Xy/sj+bIske3nfhzLgpko0TqT50X6qx9RH6gTDZfelF1Zh9jamFNVqm
qkDLyCu4HE3oBKUOd/rviwP96T8P4wIPWBhSCQEnapotFBQ+UCx0ZNbH/4L2CYtTO4yrHKY+5xB/
KYg5Hjb1kZtcyo8xjX/C7lFMXIDtq94FK/IV8LxIBq5gY9QxgjYaQTxOQn7Th3qZAXk/4d7FflhW
v0g98aTLD9KIBXNKWUDj8s16BLrgQYAsbk7TmMcY9BFEnW56vPiY9VLsjJEYMKP3BTwIKWcBHEMs
wgwlGl4T3MDwok8MnbB5J3IT2fVFCxq1ho/YhKUqXLjstvJDarFhhEKP67LIeDSmAw1uF3qJbEXB
GzeWfBhOTg+bdzSKAlOdqycYqfap9o+CybdWOiQ+6tgSZ5kNsYqNFQYIyXKI9JnfPgEj4Umkn3p9
G0drGZgig/7Gith4bDCHmKrI2/reTpa702Try9yT8UPqFRRAAnPSsu9bUFyLNK6ikpQelpIgFwEg
gyvDnI67WgancDbKkvxaZKvSsY4FooTBCB8t79/mSDDpI7E5moyUi/G+ve47FNVnL+Aw6CcwzqY+
LYleOgtpLvLOra3LeP3iDTHpjf3xP+HZBElo9ACPsJFkRkKf+BvY5++hKN2DyfJIfLorExlTT6jp
co11Rhu71cY3DR3sHvOPLHol5uy2bxcQgvt6oTfeXpa/NFO2qn9ngZec50y8WoU5Mu5wDapRFAFl
04pxX8xDLZyX+2BO+JzMXok2MWVw0CaR6vpE8fynAtnHBh5q+z3bn6ZTlpU1/ngo3tjSJdeE0tey
r7T1U3p7l3K787MuaJN4ah8odKQRZIu/fh7nIRMvoM3mcjgVFEwW2Xp0FXovLL3azVAGrUmq5QYJ
UyXlg/5TUsO2B4e22qx5TfhKGZi6+NqF/XV1CeDGWBcFZSfXO5r+6znbDXj8/2J9fW2nIIFu1vWy
y3Szxb06LNGjf+ilTaA72W00NeviYcDBv0BpkrBwGuuzhQm8FiZsp90p1c4zJXKDtBeK73mOWdsS
ZZ2sJ601IWS0qZm7o2anpM3fHn0voUBqAWpJvhsmUJwZyZVYRRaIM3yj3/c0Q1m/JogS++jBqBg6
RnoY/+uz9v76lPQa000IU4OOv3M1iv/446juIOzkqfmwlAJGLKVbcIa2tlGBBT5sYdVyUnbPFnXw
AuOfsWwUUbeC3FTcVc4E1Yms75LlgxWjpSU6PhuRyIPT7QaA/6nW2uU93n5T4vHT2Y0Gwl6EjhAZ
doJxGA6QCiSIX6aQ73NtOP/Os4qHABc1+7h4BV9e07gALpAc+Chjq2FCp4rzWEkphlEe847wxqVZ
XlXp7CRwmAdAN9bUgCJ1PQldL3e1t50wFEQkCkc/6MSsCkR4C+xpSmk3WvgSPpdBuYqdxhNhnLp2
Im8IdfbLsmyfeIme4y9T00Zy7R16rWbZqaGA63n//7sC9mnxrrOPhyRwhZ2gbAgglS4E7cozWgeh
xjkWuHaNJy1jIcGcwtVmtWAqz7N45pGfMT3hjGT1wOvKwYdfliselTQITfCGNtntgfPycUdBOGc2
aU9eBNn9tk2tZThHSveMhv9LuNXf2mNNytYUdowiYhiCkUnB6tUtYXcAMpj8/cyUEMIHPC7k86jE
/bg38j5PDyZq4FmTdtjgWvOKWBZAhloJsEC1yh8f4H68u0S1hjPe6qQTzSqfRla3Mh+fKjki6AvX
CEC3c0ggjPpab/e6ufAbN3CRYZWBput1uqJBsDzjlogsfvP3UF6i9aD5DLAEh7Z5wAcvtzG8Tu5Y
cwqjlY3e1n6Me35Lv/flZfKeYN/Q3aUXp/q/kF8kT/vtAqlFkW9CoJWK05iNkGjA9wYsvZAlq09E
xORjh+3Cl8PJNH3cmTB2HA6horqHMqwCbOAKOuOXduB7zeeazETyTPIMnLHot0ncICyyyf6bLyNd
E42Dm2ed9w3zsoReMJBo3J/H5rXoSXmH9rhe82LJyReBD3pPEnKbtniAG1xiSToXuThcH+gHIdRs
LDXlg9a3V+dkQj75e/cpP2KH6+PgTc3On8L/KC9/FrP2cNwcfbn//86xMs04KounS0DaoNB3CeET
kMwmZOyKD+QR81DezeiC7D6ujb5zhNmaFnzODb2dRZuZsdO3YyJwGM64Qg+3Agl4r28taDCEtl41
nWQSIVGYfo36v9I6uusnaEnsMaubAznHTBZ47SvHMK0rkh2UOWSo9KMOcpndBM44NAVObP9Do0rA
uGwyvrd43fXVS1bNc7dTgA1CE02ITTnWtRAZOI1zYFkGJcbu9G6Rmorg+GN6wvRSXsP39VhKiejK
FixpLc/9bPW38xnIogkSL2ck+n+aGPVL0r9pYD1aaHHROxBjprYG3mjFG2EiDqpndHUrriQViXYH
cc3dbPxmp9MOYfjVLJQjOLYCGnEWxGzgLs/ry35dofUex3twRZE5VGZAAZrixdTFo33HEme2zGiv
Yf4Agg0/mmm4YCsaazFaAHVsWMd1Ebpz0lATBRNRo2/06dX67bHG9v3ceiGzU7r213XH+qqIM/oS
t71ElMFbfZqIf0QXyomwIGGtMceH5vpWvYuMP1aqk7q7GmqBS33KM6jLLkL0IEUFqibqO02wTOe9
75kCJw0s30NebMnmSrpu2v1lDM4PRC2OF24qu8+gKpAIsHVMZdhsfwNJIIv+0Jkg2d4lIVswh7U3
syj28HfhqWAV8YD/Rd6OPFa8G0K3qubgdwTS7ff8XuepZHwFYI9uOglLnbSBAPcA/b4FUCX/9YJj
IPHPGqGsQfjVbQxT9JVGI8WwehINGMSXAy/1XgnkseQFdEGBaYByL0STNTrBFFTlpxgnlLk9clXD
8MWPbfloz5OJBQ08VXyNKatk7Fyn2q6HZd/abDA4oxnLkz0SbIPRFJIWd9z5FuYEBJsr48RljURy
XUGjTzOAnMizTkA9jXt2DXkFpXzG2hwSuiQky9uK/B5/B9pevmbya1AxPN/fjoJ0cUHA0KhUL1/j
TgJShaErWoPfrfTuQuRNjt/5SaIPqOB2oX1bhNUQN0O6ExJNphCCVKSs4P9njgvGuqT9GPr6ZkgR
UKfUoqceD6SkFi8G+PCG7afcDBs/W7WIYcrShNxUfsp3y87sNnQkshWO8noMHrGgGgoInpmrBiiy
MunVPxcE2LXYPurAl6940u01SjQ9qOqEW/So2ujy0zaNXWrLOadYBCQU/0+TlzphAxlqo9Mqa+ql
rdAI+qBjBhfldrp6Ypyw1Ltks8lMVAmbdXGdF6L78df05q9FMnUT4KTprl72Ct7FQwLOI/T3VnEA
W+DxdDL1GOKzm/pxPqPH0p/KhQsvjR+K9qLFynWkEv4kRkXYDzzKtVNMZtyUyqmrwa99iJgWWwKN
Snchws8UdyG9qdy348iioj9PuhCOKEZOVEsldEl0G1utwzQ3VYsuSVZlG0prCJYClbNo2QkjB19q
t48ZogkBAQn0qal9qsA0F4l4M3/P8N3wZaybur2c5/ylO5QQKXrDzdQQRteLjGtcJANBTctRjHfL
Ue9J05sp2rEDCmiojLOK9ch7Keov1P/MbpoOAElONZGZUDFRWLD+e3BymQ4T47STwAyFQL2KkBCx
x/sHnBKKJIzGVis6UXT2VTsuuTkjzka8kjHO30XLLxUi8lfp8ji7TPM2ejc2C8YX4tcRXaMxcpDP
LqT8NdwvE1c/bk+ZXjcGR7loP68Dzc7pKQxWORLF1bE3FN2X799dRgNw09BZftFCjAOzxASIWjD6
XPJwR+kdWUXV2RhMUINko/EwMN+WZGFR3FDWLEfVCKAUnIeFf51+CQ+BMeFagpQgjyPxp4qF8Osw
wXFwUw35BJh2lRnBip+dBSylgfMIDdzau1732X4PYlJLmDmGPdyKl32y1FB6nkmxjjOps6eKpj3l
jkrqXiMugyOHBPGoLNnIA7Ftrv/9f8Xu6lKbQ/6XxgzmaGDH7BPEAJi8+fdInavCy4F6nlVMEwYD
Ag3svcZPZneWOS/E3mLBQvizgU58bHRcR/EEzZ95gmlmSz/I/KcbDZW0WUcjyUuEBCN4wfu0iv5X
5KBHtt2bzKqfS+lGAutVdxw9DeR88zhoj4dkHe1mrTWl4NGvPkFcDNDv/5Jkh5OljeqDaKHPACtk
tCNZUlwQevYiichIedvgOqMjFKPf0kUDFn05ZRNXP/18zlQynw5BN/s2CWBU0UeRBNPGmBkUodnu
UlnGaaTVsza27RvGiO9E6sruNXwGg6oBklGuHbA0rQt2EYLKVfd71HozWnRosRrQZRMFAThCo3AJ
917boFccFcG+A8kpGdCh/GLdUJSLI+38PlA8uOUmO5yT7v8osBzMBWginSJmV8wi5/TgqXem8qB6
b61d3IotsOrFfeqXtALmaBWYhvZ500LNEcgPHL1kIsYUU/E4axTGpnK9KxLJ+NVlMdOwaCpDLezj
SaBJredvMzwc7QEz5ZBxreOt/9mGqRZO0RtAAivWDLyFJ/yogD5boROjiHV8cQV0tctv3SKBwz+w
HB1RhuqSukfSUCs1ja3JcBTwAlgSltLlkEJyhWsfnJL8plLZtJkRBt7xFYU3pYrVoSfVSNXrG165
UouULfnRZX1zQ3I4UG25qcq7ukbW1BGnSBGIF8PM86lksIdDxka1IlG8dOQLvxCzQKNKmsVdtfcy
SyqqL2MumPSbAMae5ugT+3T1egA+xvDayj8H+pgITNxfyqoWJHAXLPbKTKA9l9dASTSOp0x9+vrr
TFfTrC5ohibNL6bo8D8Wi0P/LwsTj94uPBDLt2pmGxRqx/AI+o5TE2tJeAAxlQ1MbwIZVn1jcV6y
I723i8Z7ehT2hVfuHNclQ4eb/sRm32R2b6vfQ1qKcSr5Y6jOD4PX07aqKVoolRY9+ku5YQ3pI9Nj
l8Dc6tFr2xHw9UKuoTrblPvAUPcyQktyJ+luVsu9C+xqDkiFWu8uW4y0fCOdlVf97crJtXDsXj4o
fkKtfor9uiAbVFsrgqOeKVKWUmyfQTTVUbia82j6A7vR2LkmcbSopfInrB3ypKbazPAJts3bxqlf
+oIiR7YrnhDXKyMEj1ihZWCJmI9I+pI2Xyw/1daklbfvbopTQgCPYa8o07LRfZc+LJLj2TwbUuAN
H1vZtHWV+LtWWf6N4mAfqUIWmnzRGccqaI70SF5i1USfXY0wLuddnUSWzWvfr+aZhU4UcK3vvEyM
ZWHWZC6Zv1wHxCoFQxoWQS3teQgB1KF6pkBt3ci+++NVDmUavtY9sSIN5r9trzQeo3boQpBmnhbj
Ve7JbZB893glw5dy1fjH60eyJxF88oYqQVEK5t7G6Rqa1AqZYqcgjX1hAnk9X4sTwJwhyTGoOIEw
tNd0Cv8NQBO3WqwGonfqwZxwzHQHVQDYitFqMTgPCWJtp3kPNyv+bkjF8mXzJ7ufwp1r5BnGr9k8
OxDgx0O8/HGgNG9/od0nYJfl63gJedCy328unz1WFTQ5ZcmgKxbWOZwYxJInjpXXGKBLNURL5E0t
ymMezZK4sUCLJ0oAR4qyd2ppsKf87b6EeB66lXLGwY9QsdXzrU0Wrbxu6ZM+c/IHVWuSnZr+NqnE
K7A8V+PydrtnvfkMYllyYt9PVHc3GKJ2iyGMvs3SzgeW49zr3O0BxpJ+XxmpAZzQqROT/HDkFkkB
xM333kME2y61RBLLcNrIIF12QPSClmMHZbhdTj7+hIe2C+0ZiZaqs4jwXw57QDyBIRmowVtN11Rs
yQfuWEYzYJKQ3YqC7ZvWaQkBVtuXmC1eGQuukJQPJovS/AAe9gBzWbzBhgCASR2ZHbuCakRAheKd
6QUymtahbKER1cYBZdBh5hndjl4+mXSQzw+czzWAdh1erfLYA3e10qSMntR776K1q17w5B2e3S3n
ewESZmIJ1U+Wsz2N2y6bFqfr7I8JafC1aDwDHQAxCb4n8BLexteRSOu+Z5MsT2sy8QHtOnkOMTnr
u2XAVk+pUkTaE8RiFhWiprIlFYzqq/n8WU7MUk/Bt/sabKkEvbNnmiJH1t3Efd9UP5Gp7DpApZWr
E453tqoY7e1BH0GXVXdVqtPdQ8W8wDsyC67AgMOnRiYSPSUUB28UCmxrV+olWNSWGwI9mIIXD403
6uJ9C4OlAobWHk5HcG5r0maQl9KucQqWAMVMG9GJGmpUs91/eDsKXmCoFZcKWE8khwMwpDR9KZoY
AJXF2eU6zcDdtlOtXb72vgSAfvLWPmBoKT8jnUB9m3DJOod7j3uDtjW6PZIj1tht5juU71vT2uId
nYn2d17uzuGGF6kzJV/rlat6Q6U2zOtlo883QbPS1B+TjgESHn9NpStHQ5+qepHYX+YirZJQ3Mwa
KvRSlrEpStmyY7yQM1MqP6uiZE+eLdDT5ayaWGhGlt0+egG6fUXw/KEG5/50SVET3Ddkae1yeX6u
dtMKHVP3Q8rLy0FHQMEAtNPCJZe+kLsK4QM58LxThBdGVavrz4QvsvLX74ScjNfkuZYkV0/rIQQt
95S3jtomNkSL9L5TqnxwbN1/+kovzV5paCMLPDsCaQxUn1rMvddNdrF8o0o2ftdCvNIaXAXlCwkV
nyWG3w02/1fwCZP9aQD+Ftj2LWhSous9sczkwpvAUdOzmOPu9Tg4DH0BuFKn5xWR5yzPLblyeKWj
SzpNkJiYPibkg+NbynUCJDJAo5eyJ4JBioFwhO4uPPnyuS4zbRne4JBhgvZ+tio4ER6S1sF0PjE4
CTKdDJ+q1MiBgH52MlZaCrp7ZSsIZNkhJ3vO71NKQmtHetpU/o5b/ZpHPB3sNSd1wCA9Bl2UpU7N
ftgW66RRVxCc4a1j9pUohD+HMj1GUWRHGb38NllDeDD3pbNulKEo8US6gr8b2tIOkcdgkFqxJ42H
OaUTJlFvwL/MLc51zXv69rFzlX2ekwzEoBIn7GUQPGhoGwh46yWpI8bfBSm+5DtPyRCyS1wmvRGj
SBS26TUPyh/ppfizrUQhdvcln3Q5ZZQRUB0VI46I9ANrRuYkAchErO+Xs6n6fekfqWnZRsw+hJmy
hb5Wg31cDAT0aGGNPwk8RNDgGsWeXt5LsU/LeykgRdJo1Y9FzH9CP5dxn+AN/ujj5LxhvWoyahPC
vtoLhaCk5kGMuwYmGnlisIfRDTBruDmE89DR1RUmyfOYSKNDv4zsPjmA+m/DoenNLOSHH/PU4I0v
OC7RMemYEZjZUwxM3HzO2Zhu2xXH39Y/bdJb8mQTgL5yfDl8ALlIYU4YGizhCtygpz4jNy63L/xJ
OQ3njEX+sdZ6zz1g7PoiVhJ1PJ2Q2ONMtcIBOGW15jds4QDapbq8FlkM97W+Vmrkt4cj8/CsdswG
Oyix3WrgIjShw9AXm7UZbuG2vlESFjuh8ilbqmq0+MCTAjpokKGYiK/U9btLzVhM/ixnTr9sIKiv
QV8C42KEaPGXXqimRnyRBSplR6pJOBsgBlA4IAZAYvHNkuoMPhOafUJAeGrYYXnd5GTMkkhGX4pg
Xyleyf+tZWUDoDFFO240zxz0aCCZKROwAEt17WOJKYZ2nND7qebUEBE7TsYc1Jf+k1hsWRR9IX2O
JIVgREFnsaHU76dAROCaYMlP3efuahm1XR1W+ti6QZjAvX9y96kqCbXUOOeIH9Jftk0ZYT45TjXE
KJsc6AyD8C2v0+hCQrKjA20AgCpmZPOFiH6vwEzGPBjocBciBS16qulXLBfiOwXDpt24YZ4FrWkT
jEejvoTNZfQ3X1zikaFeRnq1NWjjs/kt8VLqF1fR7FNCNFhat0mCTuM3RB7SvmgOl8K/ZZ8imw0F
Y64WJoLFleG5k0cgMPWlJAokVbKnQcqg/mWOFlW96/Ln+PRCyN6kAhMIhmP9JCF0jIGHFccZk2jz
PgrxYDu4iu4IrKT0HW/ZqWl+SB0VMsS4mc9khOLSYHC3CeH9SClH6DNDBKKnZ4y51XkfOb7uUrh4
ZRvYMyRLonh4O8iEHCUN1LRnUeNA0u73e/BFYN2JYSTSdnuJWqbs1m9K6cv3yTPgO7Xe1Qivv+XC
DCyiMSvKH9DvX11hRSIaRqW6CM1NvT0Ad2yuxlqskfFZV6rCa8BlvL2RtV+l9KWR2VjiPzORmOUY
5CVnvG2AaXeMWC0F+uwXHPAjHlzW4p7nXeDHulv4uq/ECBnrwUJbJMwP5b4wkdQgavgT7a8R6Kmt
+i7/owbTb2i2o8AsR7IptF4d6E0h1E+YatVn70ZGsxodpkr4CbgwaWuI+YtcVEsyTZ2DeIdoiGm+
sQ17XOCwb4h7nVwup9FEe0X01AubVMGH2ywvsYH3RnphnJG2Gn/XUM7qtTxZN7bmAIwGJ0h0J/xT
+5lP13aGeL+ixPa0RBA6CB2+0Z521TJMroAJ4SDiaw6td7yfz1mm98WcYTlJsdr4FbxzxmoEemrb
VYb6HkplCkykmy637dvuvLJZgBVLsjtaI5+Tpuo7m6bYTkIzkkMhxUtjkbrsFJMrqV+kq7AixgHJ
Lee6DvihLCFly6mx3xjM4IX6a8ISo3IR7GJkumCWqAgXMxJxlGfxlQDbm9BKNb9Pno0GYcT3dpHW
DPzljQ5sJ6janO5rQR/NPl+jVEusbWuW8eWDF2vspwI8R91hK4wdXWxd8sg0YHHJqWAH5aXu6YDT
l+AmYkp2UFsHx5EuDdYROdDRveX6PRmfSqTrm1FwgwVb+7556cZdqCGChKXAZVoCqhjagnoEiXSa
c0XrEHkknlR1RCtCJasb1J1uduDZ+HWc+Kvmx7h80JjFM2r2eFNrzWrS52Mf0QpViwwDJtEi6ytn
ySStHvNMf1ZUXSmKTJW61qFTCJprB8Vu2LjX5j1A0R7fC4vSUucAay05UhJrfBBPFMXqipqHMolv
ZDAJQjWkz/pptP+1rVlVIWQ/j0pheiPh87lvbU92ENOAtHhRMIE4QAAioKA5AT/ffnzAPGKfVG2R
9Gxl7aMSjv/5ncEjApWKgnXtDW4nRcpGRX0g3bipFTIhETFiRMhKA3s7OWZoHeYMA5peP2xmYeH6
Une7L1oP3QKaxsugvgeGf+I4SIfD1nO6gjJXxcMgPGiLgQxgXJH4Wt6h8Uhc8WDEsyFFXMBE8LTp
HGRnC6zStz1Q0kvipJ/lby6yc+B/0i/keI4fTZhDp4IJt+x2zwif10Q57bX0YTJWrv4xwnrz6g4e
+3I9/10Xrq8ER404RVq45elHDcLtnRDv0QfSEUSrq54Cl1RVLrsku+6XXU+Anf7buCbPXyzOBMm+
0rZK+7mtTCG4AvtuLjjEKYZiZWQLbWPkHOi1KeCniJMuq4UcODJG9gYlnzGMSCmy0GVMitNGEB70
E/Tqmgf7WlDHuIbLdoCukF5fgq9Tr1R5MVy5AHjsZz/LZlK52Hr9iHTwbAqZuSnaD+0RaQij+Dqc
GqmgjnplI3Cb1DBXNGcs7t0GVYXpyIOlLJe1FBuq4y+gAVoGNenuGmRKfS2xzCp93Eg6HagrgzzW
GryqiNLWW8wgqueznLeuKyK+IsOH1a4fR4XNFGHre/vkUpr5pMn7qzK/AnFZKw6BmUXKdYuSA8zR
+jlcJpPsfs7lQQt8pttkzk/R+EOKTAc6v1h2/gnbXD5KhX8pZ9pBW35nF5ryk4FhXwAOdJN9xNQh
aFZAYwFlIysBf7PuFDsf6NGergVdBAc8XmE7jfVcgZ2O5WgWdnsGlSsD/Yvd9/pS0Z3lCRkIBlfg
MdsSjEVEnsWnHLZxCP/0K+VU1wPTCmBBiRKsmnyxtiAWW5DoeJUL1ZdXVp1XyxH5lVeTXwb/3hVx
Ssh4mtDlWF48aiARrixeoRRwqou9SyuL2uiCwQ4SIzNU3UgM7PBkIBTi1XS05PKH+GwtJSihRfQa
GU3XcrsxvkI34ym3dFnZuaZpHBq/QrVXCXHC1mmpdj0qydUcNGL6JlB/IpzELI3KJbjVvHT/ALz7
bQkyp4+xvAIXP+Lb1DvJciOpXcEQZDnCilrlweDul2FtTeI+o728mvn+zAGdp/+26Bic4xi4cj7T
/JL5hZ7UkhBwnaUt1EMps3tGCQQUXwCJiLcZXiTaxEf7yXj8acdjRZsHF1fXHAOty/WAdd6k7B5t
W7PQNPkecOXq827PNWj9KXMEAjGIpvQsn4AfUOCJ+xgGcRqOrvMVv52Up2EGOhWSR5AYhQz9BOib
DY7GMvUcGI36X/RHCE/bAzS2UcOioy15t43njcWVYR2pYMtwxAGcGDiN8cEt/c2lKaYLRoLiDUhp
HM03ublFeVQ4S9vrgJxxfnIykpWAD3T1Sj5jIIXMoGBnU6SCfFLmeEewkQIItpO/96BZtz1Pu3eg
cUw6kT08nL9MC2Arr+Ooob3bMIB0KaVcgzwgEilVUkePPWXa14SUebuGl1fTKX47u56r9T/yOfK/
PcoSu3gmcqA1AGV6XTj5HvBP2GjtTFaUY9lJBMqA1YdmxFqntqoWw/MUgvyQ1Vv4hi7HzHBuqsei
8cWUpqItK3z1Yb3BsrH4rStdzW6EuJE9bAV0fYyDxlf6ZziGd3UJbNnn3lY5rrjzp76kudVv4+Mz
hAHdykmDlQY9AECox8dmvq8ZQCpiG9Uysn1IPkvANw5mfxFJuNDEINqSQLzpy6fleFhlVO+XAafb
zVT0gFaCxDzAwqAtDmz/DBF8PWFClEYr0jDiW/mDyJRHR3JgDi3w4j77QidRgmEqVdeZN6CwNKJJ
UlBBOAV0W+cjuu4U1ojZtPVc4QcxaHARQ8Frz5E8ps4n79P6aX9H/p3XUFuTLfyvme24DclNTW41
39tTk2BlopxkDHeYWOhKE6prP7oPo+/6cDqwu23CFo0fSOcKw+Fpjhte+UZSpXA5jlAKr5XxLuq+
zegy+q4k/MwQRpRzCDG5X9c+PcOSMV6alFtMacoHZ6StEN1P53Rkm3klmDhmC0J5Mvbel3EnWntr
r6G2mf3IUgKUN7goAWlewcFWECSsV+sHCV5SOy1YbFSpGGymCt+CwH2xVY7semzeGdyJHeBQIDrs
D9yNM15aKk173K+MNUwdv2NWs9Vblz1VEjz8LSptGjw7jqcbxIi7+ddxdT1/aCPuwvjxdzoATu8K
iVtZT0FSlTTQhThYs4B6O1uwtqRBctbnwlKuCy7FVAhocGm0SBrBGLyoTH3PA4bGP9AlIsuTqeiQ
VCtl/gIWJUT+aM6wYIOyl6Aj4HXTNCqr1YkmwmV3cFYzlMjn0G8Cc+tM8AHl3MRcEpc7Q1jpCGFL
sWLQqfY1FO9y1ug/2fW9CMDsq/tlKr8m9Xo/r+dqHCcFmHXr34hCXBlGqGa4PzqCMREmdobRbQ7I
nta7QpsC+PlcsJ/F6vZrh5RcNzucwN4shXS4RNCkaXgrfNFfOWvLdkIw7Gozmgkh/B2xgl17N8gz
xrrSXxBVOuodT2553TsAZkvw2WQooktYPkN5TrpLudxVOmJzhQZatV/LhgjyT89OFuHr+GsI3882
hxcsPPOy/vRX+JAXzR4KeE6ACY2+KePvrBkPho3gYEppob/oNQSvX59enlZOsbKe+VkobyduX/Nb
fn4ac+jIl26zvlllzelglsWTdfC8adSXtdWo5PXl9MGKS0ACKBnT8eWYhW6A1OJrOp+lEtaeV5T6
oIArbitq7EaKlcXinLGeWytHNiEdRHqLmS3x21oa1bbmIa7IRmr5qL4UVP61u/rruALo1xGTg5CX
6gho3ETw5Nk5DhWozwUl2Oe9LCBuVfl2YENkIttULOJIldPwIqs7S1SFaEcWvUN4iTJ3JGyECwVb
TGdlG316TmflgRfHTLO23VPAzuUuT3l9EK8ioYg/m4ewOqvIJVDCbwx32K4IePC5jGHWuMzyZba1
lVZ7tgV4Rbwh85yevmFTwAPLIQ8GqPJc5+oCsR89irVWQ6f0MailvBmK79cHODjFbo1oJbiC87y8
8NazlT9HjFVB+9j0F7/2nufd1gxzT9o2s8RtXqNjGQW45XjOxCnF49mmcDwLRMaozlRNB0FZixa8
5KhkrsdS9Ua5xhmlD04PKHNXqdX+nlFXJROw2x2BhsWIk12tZRFga/Eb9GTZUHUrm5wJ98weptUS
uvWEiuvfaywpPn76jJZYUzM1Yny47L7i/2BH5cZ1nwWOyN340PdG43dl0AegDY7hyqfyO3t/wN0N
E38ADpGdCVxb4QjEPXAHRGQOthqt1KYzM0xyKc8fk4pAJIfUOzV9DiXSOTEMyIU4nNY9k/ppiKoG
PQPL+9hIqne5OmxI4FeoLCXrllrGxcHPXVCHtR61OAzlytEa6ZDNA2hW7C069E889gLvUAx/ZgqI
BTJD5pJ2yc/VROVEEUC2lF6WWgXYbaiFlLdpxdTocDE5NrBFfDCQIVEJGBvhH9zzD4fXQGy08F44
RjN9rPmCeQi2/CbDOD/WwPapTi0/fAA6ARnfPrS5CV/5J/lDSWjzm/RckOLRHqs/zJhvXqx7Y+S2
vizAVPvgLI7DlELeUMUdyaGr+vXlgpUs3pCzl6xRXz+ITDJwrVv0QRT2yy4sobjT4e3+a9LTnntE
DuIZhtnym5e/3gpMeePlrGtZOYh6vTGN0WmiPlsMnwLO+nahLHKc0V6FJF3x6VQFwyaAE+Ca88G9
mTa7jXosgpcRwU03gNfSNAfsskQrLYkIvzQfRJWnAJS5FtcXNJ9b7OwAQrTOvFnTXO6G/je4FZ0j
uvLeh8QQcJso8R+EUcrU4f3hjb54tqWZy6yZZ9uPvvaDt85A1mMY/J6ZTYgOu9FrjT9Ouy2Jnack
3/LjjlzLacS09nBML+7ZSmhH7s5fdCu/rQxRgV5S8dc5cjvJRCgDr6mDVDCrNrRZ1XN/TKjJtbDg
rMLcqdjI5zBc3ps+8q3rHMEVr3+byL7YIgaij5KQpBxXfRe3mFS2wUgrb9QG/6haTSmLqlPteuRP
1sRvGrfBGz+dBluEc8AJRpo+2spqBWDO9FJ4rYWhZGwbPywkW5X3Vn32529IZ/Bm16ppEl5p0MO/
oPL0tsBnRuLfgPiRf2mSWDfP6+kz/fpx0quZdBLScAp2ejN9pBCaE4M8kI7IKZUPH7so07V12Q1M
P9tEtvvKY3YRAL5zqjLeOfywirSDMWPOvAK1VDfDVjQanKxCA8PFi8daIfDTFj6KPApQDV3pOST+
AjPWqdtOLTMuetmd5DoKw/yGyAD4r2f4yfmNRbPOEsUlj61p+LJCfa6vWYbFZRoZXmYkBoAbJvbl
ts1gbFzUZO7kkb1ooqsb5uVGF3pWf3bnHDfzgxfIIcvLCeIZassAibvL3tDZqyLSKE5AZhNxGeJN
0TvVrHcnWKHnX7ztdb1M3N97duwvV2RoGQjcfC9Fn3bF0Xe8VdhayoMULKlvN1AU6jH3p0j2f2iR
Qg8sIthv+SVs8X599eq7XZhk2OVBs2TF4Apg/dS9JwmCRsMlzJmIHrtffG5yoJsGcTtLEdmkcgHt
5TMw1jswRWIWvtJ/hw2TjLuDC41SVIOsCTcyFJMfrusJ1BmQS7oqnNsEWXQuTv8FrcoVbGw2tmgd
Rf+ugV08AAMmyT0eX2D3dS18Z04ch77+FwB2s8P93AqNCraCtDWzGwda/x+QcsbK0FYbbq68l5+v
k+p0N+DBcTA/TLVgTY5CswkOMBtEasxhj56309+OrzRcZZGzNpvthc3OtWrwrj3tqZhqT2K68ZrS
38IcePCMzp0q2yRN+clxyaztIl3ZolhkpQfrTkinWk7KU6FNwX+FtYnPEZm9SaEYhe/lEhMMpAxy
QiJy1c+WqiBJzdYyungujNwCciprsi04YUntUEB6Zg6SsYYenSFOEZKeT0zcZjx/sTXB7ODTS9VX
Ri9BhtlAGZb4knUGcDvRNXf+KwPKjQydw6NNmtgluHShJMOk/Pn2D+QQtr9ioHz5kw2cMwgJd0NW
5cHIHG/i7pGuHVvVFPvCUDSj6OrDzy7e+aJah+FNXuY4Th+IzP+VaM6cCr6lTggkX1T1yMNEadxa
wARwVauRZBMQn3UFYi07IHdpXYkOwqWAvWOOJMlgRY58kWUfhDmuO4/MDCmQGcjSjZG1mDq267Dy
U8/fnevUax0M6xplfUDX3qXpjsmDuf8ZLJWAPmjwuDsG66zwIJdijlt4eHaZcE0+wMT9YKF1j5lG
n/dcRbXmTMgETVQkk/bXsIpMKeIO9nWjUiko/Kl8wohUx66NQsDALneTTBiApWLc6kFb6h+heG10
8lvHHHtnY1w38Ff/iA5rY7C3GPujIMRm7A5s8fdQNzbYwVcIBjo2uSJ/iDwcJ13NU4Yxy7M7MXwE
TUuzTJ4cEwa73xkJk7+whBj1X1yHQbHRtaEuKQuOaQZiBZVU9mDDvz2oFt32cpYUfX8qqMROEQII
/WNoiGrj0lVAeD07auh7mgfB5rGheT4mgkQBAkrq5pRrZtAXFnu0esaPIOtf+ZO6nzNVdD4+6jZo
2ZyHXgAQ6BvnAgWfw92NFsdtJEbhYQ/uSrwihLR3OyEPSuQIdqOXqMUMzCYtzp8pa9i4esckVW0Z
9GTVDmwVJxuvjITo+w47k+LepZ2gBcetKAPTEykNiWioImIzmbhfv5tDMN1pnogV1G4TDlbw0H/E
xZLZDYLlmZJZflTNINM3MRO0qiHijSCRtecaL53WldrwK2hs8KWjxD2NxvdnOB54L5WGBicLvpfG
vLFEtQSbwnP1ySTqzuVWL/Cjy8A6zdghWowVKrizoPOqg08HU18ZQxbgb9sJN6NTDHet8Ff5u0kc
6rf5FE9LCnyxe72q4OrzlDzLXrW+9B/Z56goOZjjC1Wb+SnZG0LleLoGsD3f0QCrMGpdRm3EPnsj
VpqZ+qYglcYvCzP/LSkZkuF+RLM8ByUdm8UeNu3OXtKhj6jiM92iOMESYcu8CNUr2g53SMRdUaKL
Jj3agM/qzUwK0574HV2xxefeWIOU6aI0XZdww6uqaSU9qb63PJRSSe7xmBB7+INy6xqVqY4c6vTA
IjQteX2uNVJFdmzlR2AU+pS8DQxgviZQq8icSqOIO6zc6NiyWVxFctRL8Ee9cZSQCQ7a3M3HwMt2
XWde2r2KCO59pRrx74BR7RvIpt+hbyVBMtdcHp/TX/Qo3f3By/x+zCxLTOKz4Zoo4xDsUG8GNxCB
jrGzz3w/PvdhPLR1shDQ4lebYnDyjXbwc89BDutYHjA+GUJlp1qnaMlMcxNSdTGrEDJqhKFNqfdO
aagibZc1IUc/Z/eO1f5Hlj8ySF0tmuFap/BUluFPQFjC8YXWKR60hdHnpjlfKGJKZEsGCyf1Jib5
tzxwU5GnzesGy0IYG8Csskb2oe8PUOFwBtQMVbULiQ7ABHN+EsdI+FTwlP6xMLjG/dLIxVk3UJre
0a91RW+bBVCrmIC7yZnB1ExDvwidUG0ZICjakJc7AdgvUj6dmXA27vLJS5ZC+GedZZNgUqhETzSK
PehB0EQhaZGrGD9N3R2+5Ujxtv2BKw1jDvtr9Ybtfg8WZJ/aBvyNgtREgRi1+BTqlDStrI8EMDi/
GJ0494i8CfbfqhOYm3j+KeYg3BlwWSnVfFRuywsrC5oVvF/Sal7wyQGECnuhnoHIEgp5TDpdCrM3
+CqYz6Q+cyKGhAa+xKA3reMdqj3rpHRWJ4UwXQityCho2uIRUM80Rnn7RmkwM+S2BpryC1s3AVlS
s7KlfW0W4rdaV1DVHTyBTAOEFpobUYPKfyb8LCyy08noWchJIqD7zcN/qx4EMZSN8pNRL1N5zlf5
uR8PsjAgl7cSkjyAsnUwcUFL6F/5yeIrheltNwl8Ytch2JnLs5QvTbl5i9mmYT3+jit/a3mcRjy3
GPIC31kTzSNLZ3Fob8su/++qu/RiPBKvgVo9imBJ6BTFfjJU/rdt/XgwyjLoT67SKxHSnshXuzfP
muZ7PGL4py6qMoKz4u9yc1q/gwz68qQocxmZlhfyRuBtO+IQH5D0bAalDpnIj8v6Cy8qekVjYVS2
uNQF/S+Q4dKIIwF4jA/8ys9feaEaTQZ7HWO6MB2INMoYrJDBIpPVT7nEV3yr+x2AK9WlJ/px+tDI
sXFyYnOEMqiw4LyaRPBP6uhsHUZIIXxTGsztkaEFM0CTu6mhF5twobT6stAHSLAFXoyViBj0KY6O
8a33dqMDvMnLD7ZZWnUToKo+XyphAyfH1OfrrwehiM7wI4ApZp6CHNOZ78P7p48FxWoXPvG9Bpi7
09n6UGypOfzH0hb5T1rEb9vy+33JT2h5tgDGNvNIMLYz5klWHnugG7fWEgU8HWOqpi4h/8NhoCj/
WQXXNty2+MTicfdTOQOC2YC3Bx53yTpnptiu2sC/X/MynUGBROPymkJ4mYmUsbYVHBxtIrSMdF0l
6ws6MG2ZoZyN6dmuNNqxSfJ4US6KlC+eBjz8Z+xmSHZ/yZdA3+nq0jm1rgDPobInK5nyNQu7mWeY
ZyMDWh3hPD67/CYO9Fwi8sC3MbgkHbng+EH12LjOYhxfV6MxpoPDIYb4MwLO2YG8dRouloIJ8XGd
aWMGYLHjbUb2AiIFAidrqyMI/4dWWNrKjc0qP/Ky85BotPtRZNA7SXgpKXPVfPIJ/y2h4tp/elD1
rDlv9vHaco6+40hgPjM3BcdwC4SImoaWcwEOROa4NXjmezV8j1uGiQq69N0jmBPAHH6WugQjkK1J
GCDzzzING/5fxwt4D2/BARq7SQWHH3rC6H7++n3RHCC3fjFdC8eSHIf27JmnHFmobzHP4gh6yuFH
lL/LnuVBGI/pMxNywft6rc4rDKXEU1YCPCsftsTswyRVESxmLU8R7vZz66bPAgPMa9YvmoPeynzn
jnRyovAZxcvQXnoWJAb4rSfmrnUKP+vBjzZiwByjZidHdxjoSvHhbjMmtLxuZAyrURNj+lq/Q41Z
vOKR1ZLheZLX4b/xpZMb5D72ck4nECos//KNmj04zmCxSv24gGkrEizEX/UAk1OQHd9SHilz0Qn6
NKPON6fCC5eD4rN61+MI2YyzWbksjneUO3GS40I0VBPT3E7Twzbr9afg7p9KUyZwl7bLem9Cq0uN
fJg+NBdyyLrknxI4lkVdlI9FnJDuYJG/mYbWwFVdvgTIvrOTaR7cAZixaD669zKurTeDP7p7HOdy
8kCTBA38dzQQHDDJ3tTicjLyi5ttzYsg+BXx691t0nyo47suB+mXkJ/qr92S6Ntb/gA52lervmCL
1o1ZMALQeGx0jfVyCl2erXsVj/xOVjBLuUfwyfo7hK4oAYYSuxunL7ujemFGT5PZf+Re8+NLmxsw
84+RDTyoOK3/FQ/2lJes5dJ9Hlj61yUEQ5sMPmB/XlpnVMRwGWwjU5XQ/aYRK2orEQKANEoBWRDc
e8Th62Xa1J4+RhCqqhbRFnSjx75vGVaudEXla6BJh/Vdc1FEJHk1/YXqk4AbgPc+3snmKXv98Bsf
8oAz7GR4ULXUBGC6YOVlJisJRbMKo40E95aprGDTD9AwZD5QWNyOi3F18nx0PlNXPzocUc9ZTaSz
VvHz5LP9/lkH8xwEXpwVoeBPWar1y4fnQnNtkQe1icqhIgPJYQShGPhCgPy0nyBPG32fqdryzQ/d
6M4UDnFP7WUHko0GBFpkneDbrmP/RDoGCsa4khCM/DNDkI4qCnpYHCQ8MuDv4Zp9vYLvSm5hlsAB
Z5QFuk66HVx/7yQNNenr0QS6Rq6LreL6/LIwHCtS3F9AGDtcxXDOlR02dSqItnbhgJI17fRWhoeS
0D1h6cSn3L84yn79OFj24yZRTLFBY4IUfw961SrXaX99nckobkOK/yJanQnBjqBW5+A9QMjGkD+h
nzglDAuhctiRuPOnf0DePymJj89ZuxHHjSF1C0fb77ZcQjmOcUKjUy/4V7fA/2VzTPdNKp9WPwNL
vCDfF/dH2PHBdLX8IL0eaiL7pAejFmS2pbdGGn9hc23TBPIxg4BzQz+H8Cn2HaYVfHc3WCjfJlld
I2962bjXAxL6lMVt2uPHUmVk2TTTs1kjzPpWjhk90khA1pNZpybmlw6mg/CwGWdZxGfb1ZUYzhvA
BCzJjI7/6PR7qXC8ltfuPVGlrARlKG1GO4izQupMMwch98DcwW7gD+A1TltlQc/sETfeqXQ7/Eiy
GzgKJHuGJxLSQnJxgfjGMYhzEeiSjzgZ7ihQ5islQRtDeh93OojqiiGmqoX8kUhVuATYRQtwhRJG
0hjmJ1iOUtkbNLxaXk72/RqtSgEHhGkEMwxmddsmnIPKWN5NSJrdiHAnGrSyXUlIUDyh+zr+RQG6
r5cdoJoWeILuu7qfojdGbXO4Kg3vzLRiWAALrLZ9zReIEULzex4PDuqTU4CL8Bj8fLk1mgFzZeyk
ezfX4rBqI4kcUI+yduknga13PJFUVoAqGLgEjIqxk/y2u4PEgomF4bqRfZ3vSZwD5QjS3FtpE+vV
hCUasj14Ab6WGRhOyDP6w4xqvBYhlfaE6+9f4e8D85bj2cVJBgikY4iXJmHUaeK9GELn9yaC+9eH
Pe/KJrAnGRsWV7M5zfANjIWc/GaJtZ9rM0nDH9NJwutooJwhZKqnRMhAmR0o9oSxa+U2vrCDNB+b
gMZcs3E9d4DBT1QQboWJEP5Rs9liGYdMk4FAg/I6VzSkVKlu28zBAnxWVdYHnfKx8LzA2MIhNoQX
I0KdDhI1UpOW1bWRbrGRUfKwirmEjDu5GINZXwFI6ZLhDdhKJs8LiYKUimG5MpFzvuao1jvxGQTh
SssDvi5NSoRuUFL2c1KXox6p3auV9rslsaoWG95q5wKoNTvnkJYQkcngQ0hHTPPJXy3/VkBBHqgc
5gLpji9n9hM+tsZQPmFonNHCeQV6o3RleKVbclEEgvQsSEa51s6hqUpL87yzij3vVJ228H8ILd0k
KCrRLwBPrU5H5XdLfXAKEMUCrsAJPJQ+9GzIlAisdI0/46KZAvdvjHEx+loK1Ycfc+V8v76CdqUW
3BwtpWC/qgrtzYyMF2wnJ+Xbpj75OCmX8OPqiqbdX5o+UNi/TAUKswQ3OvJs7s7Cjim+omzunGzo
a+fGVQ3/zHF/uSRaUAsHwmnu7LMtzEGT+iemxrO/wSowqFgRyUfnpjtGq78ZJTTNkgpOA3wxx+wo
D43WB+nNXJsdSEq3Amanzi1TyX7y8FRCeOolL5B0XhBhd4MD3VlHMGKiBvYUMVctv8eTqgIudHc+
GJzuY0w21ZCuQNM087Ai01EYpYbhrmnk/ZDdHGHfdjk0uQ1qWgAmGBD1rj/ayEWVMRlLm9koNOjH
BV2dYXMq8+B+ZS24fTC6J7eRPkKa2aM4fM8q0SZ5PC+VOkd8annEgerNuNcP4EvcSN1tWArriN1J
q1qZByl8yIy5Y1mSzamBFjMCaB1ww6JBTvKoq5pOR8eFsQhgOx7iGJFCHHGDQOn+IPeAtQtBHnuR
ZGA2ewdAdLLlTqB8abpAkXTrnsvZlJV4PR+SRaLsOqYUX+RO6WzBESTDR+IfOfcSF7GK59DokdoB
huY654BI12CsJFWDlZxsG91cC9r9PUXbjP5qzZWrT7YdyPjpfGuTiiC7QK6W7aEcrMUwYZAmGrT3
8HbzuOn/W5EXiqAQtznlsrqPlX5wXSpTKYybJ/pOiu4cg9cEPon4WSID5k9NWBmkT2ZKPQXVuicv
Eyl0ElM5az2rA/8gm2viEFYI8wvO9l4sDEruD7VvMvAD1Xn6BhOENLfEn9cei+8vJGvxOpWuGWRv
ORQJIX0jr1isX9vBL6w9ciMCXymKFhxthgV221PdnL9B2vhVXrGA0reK1Iy6mVE2m/qcQWnjHpu9
gVcO+VB24ER9bBguiUTBkx1iOHdECkkA4BbrfSbl5MXLrHOrf3yGNdPSyOt03hD4xMNaT+tOUybB
s0aAIPFYNusUgI/xh/pymxnxou/otNveNQfbfSQDMQSoFjJsDwX0JU+0SOkS0m+H66OOyZZeooDW
YuDxycQjmHhVZpiIvPJYmS8YI6/VmG969hpM6gAy6mmv1r/8qNrbSFhLqewOgsQ9dketIss6CwBE
nw0xfDSUgizLCUuWsdQM1dUFIfIvMns2oj/F+hf89vMziM589YeUEeNeXRGpuAkrRKjYSt1AO4ay
4lyZkeviGEmq6TPOBE1A4cBnYcqmOkPb1LkVBJXGbXpDGCnzBdHYj1qCwE5ScmHlnRtLWrmaCVQ5
SfQEk+ZBz+BKJTIhjVjHrOtPxTic3hlJ7BvsevRyt9Nbxe9nJ49B8fTfJXo72lJ1j9yEXxwmsCgh
JNYHwgcgteQMMAonxVYDS+UA3Q+vZOU8V0PAMGRVQc91/uIKbdZobONkF4H5j+Xt87T7m8h2nUIn
9tFFyDADz4vDE40wx/ipxZ68MsjRy62PKTsZnwB0VXe7q7Isuwy7ubENZFxZnQpLynQTJXGHx60P
7Pu0tnmmlMQmfFNTFEKBgKdNNqY9Uc7nyIzWNikXFeuUWly+thaadarAz5QMbUA6SwMVTe0yq7KQ
g700T6RZDQlzqgVAR7h7uo18zDTkB1UlWU7ENi8iDpH4cdTsqvMlG4QyEOiFrNaVFm0BC8Kvsf8x
VaQ2F5a3T5apLzccuvWonmNv6HunRtu85cTezU5dPFZZKLPwSXDXkI2lYPeWUr24FXklUx6/vlXG
TVr+GZi7EbvO1RUT+gAXOhhJB6Q89qPRkjk/dqKiM8xLez89iam2daIRxGFIgLU/+BhHMS3qc5li
AkFggZVo4YcJN0lsnew9UO3YNxOs8Hl8PFVSe3wx+Mm/uHqUrLnBC7Ij/IIvzg70I0NHQ9N6UYQe
Emvol0wBNr/kxIvc1zbHScyCw6kWM1gHI/icbAHbLIIZC87jYwzrfT+MmpCtTZmPFcwq4DxRyQXR
vRGlESjP2sdW3EtxDIKrsx0qhOqxZIqXOAsLZi5lT3yyVfeC/SpuLp3uMRk0JM9pz2eYm9hntnTG
RokQWU2W+UY8a/aj2ar00VAjo9dQLRUyHqDLEkYV7ZaoQTO78QAbZd+z1cD5wc69PUhh+aeRWn9p
gWygsa1stAkQNc5IfYy92qxNnX7xVHb2loRN1ko/PTdV9BEYlDcut+Qwz2rZ6GWaBMILKsp+cPU5
2VXuLbVtf0GAwecggyrnsu/mn21JbMRqXbh6b+7qn0DEWr0D1Qgsn7eITJeGHbP9Y2TNJWnWFdr/
nvWmLmSxStu+8Qy4rMeGiNJ6dyEGqqTr7/wZ+TgsEz4LGJnQTlxFTaLDPQpWkB9be0uM308YHBgK
zf+Xgb5hvAKUdqE8BVUyH/dLw9FX7/0akKekWFv1ZyV4lA2d17d2XlFDCeLi/jS93PzzY/rToeWA
j/ORSu/c4Q1fdeyWJLcqFvbEHeBycaDQCc7uoGacJXuM7PukqezNwuJBWu8JW3DDBdHZfRAgy9bE
+rdyDpflKhTrRoEUx5i5iFpYPL3bA1trtUCjsi6484SdVRZjIS6LaJpyhlO7t7jQDlpcKRfa8006
/1wsPbS1PYJAD3b9cYjbIGRPr5OR7mSs9zTZ7V2P2ytytSzLrUf3EBgH4jSk8zUWNgVUp2COgNNE
wJyjqT7XPI/jEJZh8s7SmFIh94yPQI31iRWx6jvXLFqeCMBZgMGqBS+Yd7Q3X3D0HPYFChiwaxqp
uS5KmVCMjiQ9xerhKEO/gQ+lANIsTaGsuYAQprM2YA9iwD40SOh5ayGwcyWp72RMMYnZ6oLrdjt/
1BD43XCgSi4YZPYIsPBsRkAbYje3WlY+7qvGuxK2CwHpkXjPv9/gbVWZ7LacwzA57yR2fv+Hb3ry
X7O0YvrGGIE001EG2Tu6yqbxw9m9QHr4qssPDF3XAyRL/HJQdPcWzDj9eBsdr/fxTkh2AQxb2PtH
QTbxMSQVKWBZvmDamaBYLt3HHToXJKdocFCOJQGHZoP0ssJ0z6EBGmHeCsbl7Y3z5Kf+xo3UCmNv
aVeJO2cSNz3Q8rXaK2IJyULKZa/VU6DiPj2iQv7iZFYGa9OvO3EpZCHshi6QuXhiDPm4xGdUYv2S
N1c3v9OilgS7Xe7NkhINNwIMZkQTtGcupDpxsHVTeV9BpieawKVCq5KeF8Xu/KaKBBgrl2e0DvNF
jgrNr0Oa0jUty+G402QD/fMIwkIcp+J5Hqcl5tnGpfNGNgfClgj5cN5GVMV0pLvminc5PEz4UlNI
jRKoTuyKDOJmvxOs84I4d6AZ7YctxInRnoCrBqz1HUgcjyyTjB3Cv7yFFysbGwRBFkxGsDXrmN2I
xbuX5gsaCmWs0nfb0anWhuiCVVgCBUNnhR8DqN2q1MIDwXIjtIdObM1EzRp9JWWcenI06tX+ipgJ
M1vzuqbqOQCxWEtAVJJC0t5z5yr2CGndixVq2ej4qFNtz9sBJoebjRNll6eSAYJTorgA1VvEPQf0
hy0K9RTPwatihrxVWKPQng1jFG+PpcmhA5Md1slE1kiNIdDaVFgWdERsgb3GYJVStE5HeCx80QBh
zmB8fQccWWDpHkgOjwU/UMgMyPcAAir4/7F8PRonEPAUjf2HHbDF9/q+lDkVpVX59I/PEJL8qgPe
NW7TpWWIHQo1tLsJYnCsOg2sHV5i41j6fLDf81HoR9EmWkSANkeQBywDM6H1Ys8pIoLh2wurZjTI
ciulCEofkOMn4W34CWArGq76xX2A9lYWsrjoZjKMjLWje5H+Oi8OK8HtEcVkRxq+wC7oQe2wMQy7
4IECZiEhTyJov4Wm+P/zjtmkZx00LXmNqbcpjfTVD/f5YjVQ+v4TpaeCRZ10YRL9YoNZljSrYPLY
PhzMgPYRedokAhvKAonscw73i2XXU7YR9xdTXQi8qfmcOdzETuE0GI+NPJ/E6geRs8fvQHEVYhjG
rH9DHxEPW3FhMieX8R0fEyiUXvug3uUEm91O92lmcHyzVF7J9gSE8BKCZwFg2FQQ090yHtl/0rm0
rG3nD5/Iu9NslexLojVDOf04Kal0SRV3pNNkJHYUQeRC41tk2/RJSmmJIjeid3XN6pdnglsaS++K
ax+PV6R0s4grHm9iv5vpye4N2C3QiohduOymnfnO8taKsgwe4vCd56/Oryd+nSfe5s9RMd8WgYS3
xlt+BgQsOy5I3A01qNXMg3cq+9ltCRIyibN9KLWvCvH2fYsJ1USgHAEhXNdg7+a1sqGCfegFjXWW
We75vyi7hgaxCDjrd8pXwrPu3JnHLZdVw+ccAEBMeCQdBBCc1HRE+1gOeUxeWUQsstClqmxZ6e48
ICadTT8/CjxegTx7Ddo6/OOf5l/ZC2w5wFYtBweiqNyucjvttVnCLk4hCNHg7mtExPYlrF4SKJMP
8WH4z4RSXyRWZH/2FrLcv9fcjFMKRegELAm356PCpIMaIZuDQfUoGquVhVtJsp2ARJZl1eKkbue6
ZroVfTH+jAe1O9jZQcVpN+MfJeQA38mHkHc24sQIKRkJIfn/XmLJNim69j1uuiaFpYIZpsn1RPp/
WfOtJim0/gcW/+ZzSg/vqP6cTUeb4GiY66fENgOmr1zZZL+SiK30UJMoTNs/cF1zbPu5x94oX8qT
fmpj4XmpD+horRUoZQg8bZKYivtcI5jIWEkuiMxKhCBk5qqZw7NDdGPecSdbGFJEyJQ1jqLGRC9f
DmIj3jOh0POHmCBfCmh7TU9Sl0q39BIdybag974GGfru46v/XHf9txNEcXaiU9vNWiEmK6br4l6L
hQBrege9cu3fFSHnR1CaqG0OPQcvY6Q5ilXGqbQzUhz9daj28LKgqghzS6qqgkWs5+WgBwXccAaP
coSL88cPB/NInDfaiKxc6MnYTicCV3JaSaGdyLI3goBrZ1cMuzwRet9LO0OHzgLCCUqLDkhMfles
SKwg6uty+F6+yjdvNO++L0P+bGqayVqSwu9dCnhRMBgHMGGwmUgqg/NEAF0zPa3mpWVFSu4FyV1u
MCCAGaz2uroS5yuBtIyhfOlBgczm3sscKIOm08gnFjf04dr6etR3ZES4uENhd6AMXC8+CdHKhcwz
B8COsCrgSnWqC/6+K2rukM3l64f8eB3V8i0wD0EklxByBw/tONZfIVMwtzOcn7tVFrwhVsmeJI7I
AJOq4gJrTZTTOXS2snPrU9R1008mug/xzTTAhLYGesKI9P+wClzvGVzlRP31DXbQfH9M8PthSJkG
nFbQ93vXownpfscVcSFY6RflXjTp4jRhZ6qDrlTbYbpZsl1b0uy2vLVYLkopPyJPMagU0GbBqKb7
JnAhXs+d/+DkblR5FnBfetejLt8cFrFjbErMb3yoXihvMST5pra7RBUQV3pnyYTQuiybpiASCals
cTAjS1Vl3Xrk+Ua6gx2z6oJMS2ljZmm54DkZsDrP5LcDboqKIXWbSfXr1DXHrgWZXLnHI7cMUOAy
GqqAT+EKIICwUupVX/YBcjI+FvaRWqlsKT9dMecHicNDFa1KLIuy5bJt2uUfbJGBrGoTILW5s/wY
E7ph3HZrjb8DzZuC1Wv5WeACL4DyAqKzmrYne86ACuztKehQXeGDa21owhsSZbE7Kf8RyQ4/ub+g
Pai2hg4LVTyrq/ozfSjiw9RWq/JL+v5qKx2jvzugZF4e99Fh1jpJaZK+K4rCGiEmLVUh5EoZOEII
IICvwRPJM2kyP8kMbMVYuiKHyXaxB00kuwVNJaVEml28qGI7ITQNdTZMqJGsFiZMoV4qeEku6cxT
u3yOe4IUjvERwLeQbE5ke8F9P4dOlAcgMR+4EqBpDcasBD9WNA1aeaMZRUQFDImfMJM9Sgx2UvIC
V4vLzxiUzZ/mDopAioiB08B4ixR1FzFi7FjxBkPP6lKMkf9+vhf+7eZv8q94mYIsU0XW2HNORRKU
RJ7eh+bNGEDuVBylK+TMEyDqVbXaUszChgWI/RjKE9053ASgNlt7RPwnTY7q/QkMW4zIPsMDp6kN
7Ej5Nt5giJlrlPKXdeDDKgoLNdO/55c5TSnqBT6J5n+vLXA0HCLduY4pcrvDWUt80YyCw5y4LlPy
7p4s02dmQpJjhMbBmx7NuEwJy1umH65Hk5HFvH1LdMu3IcnG2GXMQkfPFQqe9Zye9qop2Axfcpl6
/iN9qBm8BCRXcBZ/9LFjaWSPo2mGxi05FptdHdAoAOpBdFKqI3spSUFVCxv+aK0A1eLynujCfHct
8pa6y0Mzl5amMMMDro8uhDScBZtu8vQ4J524cLA1BloMYB5qgegVpjmYEvU1I5Lwo82uHdhwrT/J
VR2Hti0NUMqTPaAjztV5GNCTVhCkv56Ji9PhKXVobgHdJs0EidKrHUHxacxxX5jHdlxvzJDuG3lG
+9UGnlJRaUVH3FXxLbF1iEdtrqw7pPwaw8XBzbhgmhUv4Bu3Ot2fDcJfvEF4O6z3UW3WW0LzGQGR
AJOFT/qoEeybksFfUX+Fpi0atWwAgB1hVD7z+qUqGm6k+VHLD3AHeq7MX0zW9U7XoT+dwePqJJaf
cimE1Modhb/nT0Ws0fJfJkL5/42qlqGgKE9s4xGylNl/d4nSDvGfgActpwsCgtB8fUw2B15SI0qK
xRq+NEpjY9ogPA2nDGCbaCQMabAJI8ObgsRc0LzuXWN8cDdA+Ega0pJUZ07gssVGPkkZRFMLKb4L
N/4AhHcGn7ZIOGTGxZDLgRX1FW9/fdz6wRDEu/+Qn8pfw98+8iAlBk+3YIVFK3MupQASJHmwVtyR
ItiHYTABDtXDfg6KjjCXu8hmpLHanS/OR/c3y3zb22arieRYmlrv/BVdjaLukRw64O4+kHJ86tFw
V59C6Zap1K8k90ELkt3R8840vFmNYfKCryOyA3ARnjir+HxmIHFKQQ05/XvoX8CJoIXNsZX8kL/c
3+KWyZP+xflo/rfdxBCB4+JEx3ZsbMJ8VeImg+mwwk+ZFpFh6aff6qOZp8nAwFIgOqdJtpnH3myI
Lfvcb6MNaNzvKW72eDmkkBo2ekRVZoAVjYVKVZokt+Ji43hMi/s22BjqjHXqzrgLKQl+VGMpn7Ok
GNp79wi0Qf4YUBOF93qxxT4KGF2ZPtdijldb3HlZ7QfwdflYyPky/NxZhaclDY3IxtQewZAGElmM
7i8Q47z5MTtKBsTnAx0jXTOBS2YrUNi1PSDXh6aSZii6nAgdecLa4gYAWPv+RoAV/o8SDEYPmsw7
2NDLRbbNddVNgwu9WBx6Yu8gXpThwnIdZszVvSNmx3LKb8xSIjM0RH33H4jXG1fDHtGag44EpK+q
51tGwdVkJU8kpNipfVuh0VaLIsckVV0a5rDIBaAblG40LsB0Rr6aZ1Nel1u0VdVTX/P8Le0EgW5L
5EojoIDG9an/nlu2FYEU3ffokhcfPJk4EJC9HsAUftB4KNo4rC5jHmZZakwt7pczle/wjNw3VxgS
Cx2hVx99GHcAtBQq03lVRtLdtWWXsy1VdaFVW6PEigWAke8wn+HHkcFoYIA7r2nrvw+Amk+MB4x/
q+vxZnxI6IaxNZasSxejR09HNSb4QJE95IuJJ8T1F79SsQ5aSrRK687loWypeDdVM6JtxQ72bgti
zueRTljiTveJqeRy/4ibVJOFKWrdm/uHJ3jbiBC5D0euSvVX454HLd0+hO2ZgD740nZnoTa+az9r
BsD9LTlk3BT7UNnmk6z0tik4Te2IRQbqt2MIHSRGGc3mh7vw8Z3LliFMCIiMVKPJ8517/qNTGBCa
YY9hXD3iGM0iIIjqbaOVbcXs+CRNJaOqYGkUxFG35xfA0wMKzYZLBR5E9hCRhEBb7Fs6lI+rIvT3
qeJc4sPiFATzVWYE5hU77DAKnw/LcgrYhgU13mWqxgOQk5VFg+api2uTOoGhMQcKYkMHyv9If8Cn
eW7jrsx6e7+/3QNeSrXXBH3CrwcuBZ/NBRfQujmZlaDCHgFX1aWpjSLhi7c2op4hnoocr9VrJqEe
GuD4Y64FIlEseMigiRoo5cwvEf8zDKL12Qa5QH2W424iS7ExkyhinM5+9e661xtscNH6c6RdyaUp
R+cl7GCtb+Z5zPn8cwjf7/XEZtt589u69454FAFH8gHESTQbKStnpk5fgwysL43nFo00fMv4aiFL
9kyeiNupH02JUyAoLBQw5G185GnBzq/hdBUrrCFUnY1FN+Prk2YcvlSt4jc/QWM+kVdDKYHKvAN9
2AOjGLdWSYEy56N2zm9gBg+00I9SiC9Kv7M0sn+H2UPcKgX4L4PN9w3PKtLupR89AuTb1RPQJSHj
7nKs3+jByOQGPgD+6/s960k4OMt9Q53Mc4l0N/24F9vVxr48sdBFF0ai5jOokezWhvDNuUTyG+75
9wwx2fNv//WcTx+qpJgtWjK92nIYL0R+poDr0qyQw3r9RUy6/SSxnMaRUuZYaBW26eVS0zX5BlVE
Q6LmAUaXOThPFbwnG+r2UNLBeAF96aHnDCb/BiHP7JJXEgpQGJIcbgUlgiTGObrpk4ufiopJdm8l
2yne0Y93E6atENj35cJ4FWVp4aOJwCamwPU1LqP+zfjx5sHBBxaq5/4qJw3LJxz4aI75WVxLf5aH
VcOQUKnH+aoQGxF/3CUZSaY3BJeHisEayd+Ccv+UaD607t6cwfnyqu2iYVVmXKCNEOvC6VzyAwkU
OdSSXCOiiSEG1QucnZEarQFQkI2H6izjaQ/WVOoDNPH1/JBzAgQTSR8snanrIvBGiZoIcH+PLKQn
RudJBCzHs8ALdirxllcCe6ninw1HBczMQqhrQ83gArwjxn3/xI66I7KzNFmjb2eg5J4DEQwFZIW7
zu++eMLM64tOVuurrIrupxgg43QnDr1bd1nDaVPEryDqwQ4j5pGRQc2opseVXtQbJeOmiL+dASxM
ZQbu24kF26UkWnRr9Ofkv8yYfsndOlXPz653soWTmSwqpCjYYemxateigfkX7eSQgg55syDXkdOD
+0XUCJzfoYahsJdv4ip9O2kdiCHlYWo/R6Wd7n3heAZ/7WfcKiBH3TNDR5+sQOCY1KQqr2jKWvnF
ezkJh8qPmIS7w040g9UGFtaniRvwV0SjHR1cJ5oWTTJ4i/8kc9UvjoW2eM6iCheIfeIYLByHfbx6
A3f8CtYVqJei2i0210qgo5k4MH58YbZ1jysYwOi0LbZktZ8aVBHU1UJWKE/pETET1kn+aeM5ykcX
P3+SZW1Lizi9FKJbAYgggQgiSn0kI5rf3qvZ3FrohmpUG14JfFGlSMmC6XB4kFP48zwIcQGv41re
HV0AkKi5iNVnj8OJ5pWSm9ikzk9mJwCJLRAGqNkY+HZzP0OoGHlMt0djn/jX0KIpFgdt2irvgALD
yXoJIgAP1yI9H8l1WdATy6le5TMgonkar0dB33ut0c2k9lpSybs7VR5odx4bcdypWAuDM+ZPWd0e
xlwkDK4gxvbliLO4PDspVKxjMAo/DtjZerBmyhoMzPR2UFYi8mvGFfqeWPk2UvZUUUedyJ0GgOCs
0vclzBZ987nsYLqoPVofE9yHyQsHvcqC8To7XABzYX31asDg3Y4Ia0tfCMHTBKYM5r48m2wxFo4e
P9h/8vdtfA0wNwM4uaRgJxaLGola/i+4nwXSayf3UFVsx2A3f9iEeiGNTWxcqM9Ri3Iyobv7YMZ7
PbS4YzPd16ZpWCFm51FtfPl2wrJ7i5ENaSbHkw7nOsaRCIq/QzAaWfiDIN/cm+/8kJM+2s3yd65G
lUEahpwxRFGZJd7d1b02WsQ8kNJpcN4R81Aet5IIUc/IK34epUz5ZJf2y+rVOFnky5nSK17nGMVW
8jxA1+ub0gg7VcRe7207GsY8QS0mD2hEFO9Q6HUtdJIJbHo4jnmeflSo0deJnabJNjiPcL0zpwec
GXzKbedw4Q9hhulM6dn/HioQRg7ZRa1qpmbcxHREhiuvTXisFqFYaSbiJ2l9fZu5HJRnv1gwezqQ
XM0uYohBInLLYILAg8BRCHFsCnffkWBcr8Ua86ornPVnnXZPFJ8umHCpVtp1THRZNvpOmcI/WCRr
htPznCZdXeqqiNcNrITG391rbBkEiNScRedB/k5pu99+oNPtI19ZOEdEUVhln3R9xOtqcKy0l9Bb
KP4nUo2T+7caY5mMV3lvdINEiZ+bTrY34AS8/E+Urwv6+vA4AkUw28OOn6zzuniMBXCX9Itbsxjq
5dOPvjvCcDchGQiPWByswLUIJOhR7FRSsGvnf07D015eIyRa5GqhPNj5fUNpJNe1gyIo1fGDTfaF
sDhiW0IcXaUajrK20YcP5WLpDnMhBjvguJPrC95mjmwSUVLhJWyk8+dMBLkd9Vkty1KTIgxhSNQI
okrnSdXgSBV+uZKijl6RUG9JA36th+E5zZLkNjW8+RThJRxOGI1WLHiAyYu+Bdtw1pLrz8aEmeF9
a294jL9bptEpM+McxldBpUNqUAzrYd2JcrOM/U8DxCXc8Xa9sD9lVb5K3sO0G2D0ZBj4NEscfpqb
8/lUHk64eil1X3xIBlqUiE3x0fixCwl7JEojsnrZSZYfrGAEAxsq4SkjwR27eVTMmcub0qmKB+0o
27S+jY5PhdN1weNQjmxN1/bVEOxAq5EA2uHdGpCqV5jdghMDcUYKkrJkOyOZU0lwzJYFC5OBdEne
3ESx89sgPLKzdr0mp+vryWqsWBV1+vmsXPH0oxUxYOiphetGyNWBJ+MQoP+VhPgXuqfxXv5is9AQ
sqlIdNkSaOeNmBPCYNhKWNeQ1HBgQKvtCbIPVYu3axTPPvQzIF1g00U/Tzdy45CXBHnCIs3LkVfz
PwgDBLjyXmP4rw3zKDnFQtz1qkXNJ87ImUlJX4zBekhl3evur4Fff0Td8XhXtSU7K7+BnCTW2FxM
eXh6thxX4b25uKOpQgYrP/pk5hMnhsBxFSdHpI2eUMLdcJg0OMhs681huXjDlIlIcqhnOLY5Z0uw
oHH/G+nXu2Txo/IKgMpaxrYJd+/zTLhxqSE05VlO3xVcj1G7jbYLsY3zGscv9OMVhSGWsiw+27W/
ZrgnEzBKMi3LOwjROwX/5zeRcJED48n4ZF/1o7a3rbcMu+7voWHkAnMQQw8njGQCSzKjDGvmzSFi
q49c61MQAce0nwnFFoegOcqthZWtDwoQXcD/0daMXUA8DXd69VyhzwKHLwI595VQKqqUAKcDUn7w
ci+bN+cGisvoGMM6WF9D4CJSPIS82FLhnR1P0B+lMbpTtVBACHTbepVEIDfwaeZiirS492dN9FiM
xrp2GahLR2M7wKwiPNoCALFNmw3XErSm4byZgA56LtQBeXio2w3u0/WyZ72asNDmou2glkOnMqDI
M816QUSm+gMyPdAi9g8esgNKoGAilwNx9kKQfECZFmSNfnfLTLWJ3hKtOXCpr50qMCq2fhmbQSU3
dBqjcmEQKp2WsTGuGKDZXFp6VZLPQvUZe5aQXBHN/xYqnVF+WW1RmDs2BEdt+f/GnxupZa81tbRy
k/xHnqqZuh/6G4ZCkTuqAv7R+XBnAhTc49wGUUG+vIXzDr6/lh+pz3saoAktw3yAfEKKVik1mYEb
aqvCdrHl+hqh6z/2I7tj9cHiwbG3PK/jK0eizKACvXMt7veMjmJdL4hMVQ73RhmpPTCu5JRThHyr
xtet03kspI9l0JjBIY4Lvu10VyulFvn6YHtpzJ3rWPxdnyO7Bu/Acl/yNWxR8XaOti4P77bfcjMf
soyGFRin3Ip+O4U1t5tOuDfGTucIi1V1nZ+lHjV9zhTaitoN8q2xCLSyyEH4eYb1eAxf17WA+n8G
8FdcZ2aK1b8tyXIe0rnRg130y+UDudsEgmmKLZWlNOXUpLtyatlCnTiFavnJ5RCdLhturb8TppiN
svqaa5w0NYuKMbooev3SO6+QtzedhF1Nay/dQ59g4mwDk7vQCVDf9BDyAlBH1JET2mREhn3pnTgq
IpVHxpN0VCRBizP13JiE+ih01Ls1+j2jkBGeM9jSFy8RlU4bno7yQptJAvI5J969CZf0VszGWQ8f
kk7g3z2PW5vAN6pAzuvi1jehJkCDIrfQ0u8ZSXZx7W+w2JjRVHFWCOOvyud1m1lVXcsTF7xWg8BP
rGsWiebkq2DtFfx8pw5ThcqzEOeCHkR4TAQAkMD5hufLAxevPGFB3xn2r407FO5aEFYLDHHoxXof
Sg6D9DZcPAdKa2XWa+NzuJQHw1mfYZs3B1VjgTl2SJRZNfNK6H0LIsz9LELixRHKBzZjKtuB+fQz
zB+F1EdzOmarrqTU/9H4nLehf/vrmisDPb6Fo410TFfoqBXuTSBXZG7c4tjvfZVC+wj7RgIme1eX
lZKDFhyFD5nKUEg8okJegRygGU7nh9wN133SahzNbzi9m6e6eNdR9TDBOJCMEoKzfACKOqKNDfXB
Xf1USYFGjj222+KV62+smHQzkXNGIXVAfUmTBJZW+ZAbqx4jo5tKJ5itdYBC6UvAQyNO/yEFGi93
mP2CCvpz2oKYYTs7cLtxnxUFcum9KT4QoIc3v0Vh5Hu7ZnEJsihTH+OeAKt5PPyBKTM9oNaIX3q/
bhPs/t5wnnvfgglF7cjQCDYkc69LcYPFJI9he11fEgLkFZag6Rc2qs+k5SC0ti4GHzm9n6CrO6/i
UcVIno3rQ+53pOIraOEipoCXBWv+RSGnGHYLCHNui3ck8mwkpspyQkEfzsayL2/bBPPKPEV0qJKC
jdekpvzCDeOaF2FhCeqytGzazCtj0NfZ3tKes++AHayHTdYSDLx7R7aT5oM4idL+QUU0gZvVMAS2
N/tPMs+D5y+ozbwPevKfpv9MxUG5g1yxy3soQea802XUfh3dlKTJ4Vvnl2wCngsAEMyYFcL+pCdO
8r2Pf6opMAbaMBBHGI4h1+11sGlGB+Cc/aHSqv+kX9XHIoO5DbUo/sJP2WF5VzoWdukr4YTd3aJl
nVaD3nV4pd698FEKb5H7qrAutv0FzLie5xj8OeD1w9lI+p9q4WZAe1E/Lg8ahtzwTTBIv9eKRkG5
B3PHAIAgHrj+RboquXdrVnsBXto3bU5n2IfdnRoO64pc8re76rfuG/juykAkDEbW6iujih7oPV3F
FMZ3Lc+zEpJNiBOeD4FHJwUXzYlryKd6FX8o6omezGG1Q5RkUSCUQbRXAmuTQezX9481TGMa2q6S
tT5yvycFAT2DcZyu1BpiIrJ+a62cJZSCjgmCDXAQeekitoy3G7uq2NN1Is9cgrLyahuEYHTsi09x
SI7c4qx25g9LxDwPe8qbQk77TCk7nobdOPaqVCTDL41a0DODxjCwP+bnj2978S2z+VT/O2B9y+g6
WEKemHc0aNdXSK+VxQmgLaiZrOSrSc1aJ9EMJtCYj4XgPDc58WrSDCVaL78YkAFdoUZ33pzhPFTX
I3mN1XA9kXCvpYzyb3DBk44eaRrIluloCTtARwpwngwp6EMIzdDcWSCiSyrkzj/YpI4NtHJZIn9u
Pn6yOIYaMwJtSh1eUnoNcHpXTfiVjnDuvIcUX2NndqA1l+Jwi85447CyZWLAFC4q3qiF7mOZm3Ta
R3wgLlCMFDe9gtczlXjV+IMmcwzuikOP+La76VNBa1KDs+KabmtzDPM8yn1+O/v/BBBvC0untVOD
4OFcY1wJRYA24DKeHsZa17CJBhjZL7zKrbzYOO6RdzXrLFVxKL45nZ/f9ZF1vXK34CGsxfvDVdh/
CxjPu6Bztzt0Tlk6uAmPgguKy3TO0StLdtXviIvMnlWQHJ1r9XB2fzbRUEQ12dT5pDZa9P1avY7n
Zmjrw7sG20Xcf0UPv0jsGZdhjIPfE1J82NVr1IasRg1JvWe6jQDncSfRqoOYtbSc9q5jx2L53UMO
GAtEkoAWiWi8wNIUgAzGVbFuI5dgBX/a6PjONZuB47KrXYDfoRa7JTMSyh+XRHMLj//Uw/IZ7n0g
9xAOvRX9FNA99Cqkq0jU3HHgXNdd7l40eN2Wj+7BQWiqQjhHFyDbHsOGHTwU0Jkl3VvmksAZZ/N+
Z/8bW6Rt8OW1iHDjuUW4yA+HonXKpdo7lKMzXlmqPyeVPO1O+o6cOJGJcahuUCC3LcI2Nglrp9iP
fg3Ve3VbGpti0+wnqaulAOiEwKMIW8e3kyT0+/UJIehs0lKlTOxkf8hygMqakAGG1thoEoUpvWt/
zSAnzg+XamSgq6TFjgPFzGn4kR75s5DeF6/GZTgeSZwSL8CYmXREkzm0O/vL8+Pd8mA9xYqpOvM6
deCzSE9UXzk2xfAtdl1hcxnyx6nwqKFF0voV4acdvYBv9DWCOL8FtiFuOPFjX+vHNeRhgHYpAdtQ
bxEA0UvoIk1JMB0wZQCTxf1zs+3u0MvPm7SD7SeXFs+ILH4bKKjbs8z0JGGuWqxppR39OFZnpBDh
2jrUjcKnmuH0x5MFBxWMdvGywJh+qRIVTdaT7z7BB0hWEzov+k6obr+eztXVSf/XZh0QpFRVdoMA
hym54sDMrSVNjVXS0QEfbjwQuglJqRCLH0uFB//y2ABUh/e8F6vQjOnZAJ4b3wwSyQmixSZXZTQX
nMZw77jcs5iXEjNjfWr082s69gVtJry83m99ELxLm3i1Yra516HPd4pIWqMYQ6SbF0AKt1+nUW2h
JTx6Xc9iARyPDJFh83cki37Tjels3/eWgEgaxxSCTQX7o5RybTe4Eb2ab5f01HkgK/tjzCM7jyOQ
zfws4M+NnkfNyNP0cp144byDc3RqoCKhhXFZqsJXajRrNFdI7kpQxOI+nvbRh+guAnPMMIOlFzsa
oRSZWKkOQf+/U6d4Vrlz33MFRRfDxqPBDH/1Rcsc4X0HaxlmdVuo7FOBkEETQUsbhsV/5L4+FQRr
z/zZpVJkfHZm8QVa7ADeaIXWmgEMUDtQwz9Yf4J8+pEa72iZSfruPUnBX9OuaLKlIOUf44bXVm5G
QYLl/E9WGLb459orx3MAIrO9w+jgCw+Ld5ynmtxlq0+1RUlkf0jj4eB5UfYK7Vzy2dRNmOhdOlSD
jnLStyx1iy445H2DDU0JFRMVwE5mw8ZlpZkF+O6+rwF7rGeCb5vvsEacUjMIW3I9LWL6J8zgIB1y
3CUxqYiQnHs/VzH5Y8GSVz5Q2u6kaTB9cfZZo2gwrqqcojGjfCSmTqkP9KcxdWyIlQJLbENOXQJ0
hUX7joWxD5xgxE9nmoN+Cz9SO2RQc9vsP3/DRJEbjM6VvXFe5u6kDDwNXdaBFRkNjG8HnhUGN19q
b6XYbzAEtnxt6lonUpk2kJze8Ir/g4G6GBZU3yGsaFHB4rHxb979M4ZFFRQ5BXLYFlx/W2n9aZV1
JaSMfolNRMY3/iTMy4jOa1zlUYICLIPlLn7ZX8SgudgyDWi5t/Qvy6HAefKFHCqi4PCC/8tGHEyn
3ANNwb2S4W4z4QHQnZRon8fdcvCwVbXf/S5BtZq/yjoWOUPldPmezp0Le3sZBRCTCWKJPy8AL3IV
2zrPee+4zC0pCtT+ZIMzqvG3HPCjYmibw8STdA/pYXKa/nmIV8/L6ff9U9FHXyflFw6xa3UEZDEQ
zvVmns/bkGvno8cpVA6dXffSVyoRrMqWaizD9lDK1VyXaAjARbD0yGdhgEkHEniUv62ArtNNXjsa
/OSaYqgEE2hRkBOKRjSf9DnfTCf8QFARLt0PQ6kydKjHgRH8IlyC6grE7ayBZ1ag+T9Fcaj7krlh
RoXpyKDlBrFuCDxT9LuE10ZnGgPiMV3dm8NcEcWVxxgx6vIbGpaR2/5Dg3McNpZP81PgearLfg6Z
JvScmTvcHrRMm7iYvbQa9pxoaV+VapQD0ZIW144hDbJWYIjEHls/2d/A2t+MblFMGSqUIiX2uJ9T
/Ht0x4QACAnISQnTsSWcglF/UqEMG0vZJLR/pptoX0lL+qHXU+M5jm/RALGrS8rwsH4nqHBl0BYn
DmB0w88ogtcRavJbBb8F3klPCzzDbUezUXwVRO/fPburtk2M22JxunqlMNYgxY+1sNRKnvkV1FK9
3wqmdRyo0zuTyysOeRp7MpkZq+EMP4q4A53bV4U3+RZge7YhnNois5Tir9VT1jScETRLf/+mDzza
g9yMS2POUBJE82/HcRQRHUvLR5MTDUoq5ARAQ26/lRsk/WdJHV3lA4x/iVg9dD/hB7u7M8YezHLM
smUkw4nh6OAD7IV85Br0KXD8iVtyy1NWQakfKTQl0wclfIn7mJ3zzIp1UPbbidyX7NxDjbTz4r76
32iYvp2WHclo8GdKyH79SvU3qULJOwJvclFI32K6YG12OssyYHvLhGK398VBlLwWE8CoyzN671+Z
8sGA/hp2tD9l9LbPTxzegQ9+S1iBG7ioU9JEvXUf5/mTBudl4zfCBiqwfsidhrmbvY4+YxT89Ej4
Sh8tDhoMLXmC+AcJ6ZvWFtzyZNNLR1kFFpRpDTZdSzx55dBEPYO6Afhbd5tv956y1mJzsnKKXVdI
iAuJj7FPHNMZ64IqG6DN6U5PFEWPMMIqex57+rET87ZvsE0IjJh2hR1CjrNTO8kZHlDVHKFCIqwi
y8ymO87qa1y9/yZCyvK7JgjdVKj0Ve+lepczsrgl+e0A/iOf/+RyGnvwA9FuaVWOOPeIhy3qU+2v
ijtX4W5Wvmyso/Q6RDc0OutDouunmAKhxf0ika6xr0inD3ZjGksvQ+wDRJ1lJQ4ZCqrJC7RBGTlm
8Bc7WujW9gDuK+eN8AGeWjv5aVsw2hFyB2UGJTn00SMuZjXPmlyxuwiF1FAASK/j6b8VRV/Dq5eq
dEhWQk1bA7A1wdAlpFxz99El2yuim/UnXBOmm0bBbpVg77sIbo71KLZYGEty3zx1GAcSmYbFZpEb
btbZ/8MZJEC5B8Xj6fo8qM7BKC4sNpedHp9a1Xu4CTB9zT/pVxII0qjGiwgAuKAecHlS0aQZW3t6
yM12mVgMaRF/dLTEQsqcViVWNKjtyCWfvT4CuMrQ1+cdIfT/9Z5owUl5V0CMZi7z8QBDFq9CD7E9
P3+B4fb48Tid1qEPQdDECRmbiKygfy4LEh64BWLdgsR8sTLFzYd0ZjIWqc4QBxbo5iaka6/EAfh7
UVa0U51e6CeFo9VenRWctNaktnGYz3AdZ4m+aWVf7X8E90hR4vTvVa4ySidaw1XyuXmm/yintWf4
tozn8lKOhNefYfpxKyLJQDIbGhpg//X/ckXaThHBRIo3+1vb+OSFOgJ7oxucx49v9SPUlj31Fn9R
ySqcPTp52xd2tHu/nXN14OAXoLG0bhxCxifmxL6hXv0EX1VmNpf21yHvQQsfD8cIqxNG4DrHxMqA
i2UTCnpiXCVg0uN1ObB31w0Vj3TT+iMsIaO4i29CLtydWrstTPAJuv88FnmbOIYfJYq9rPwLgPD1
Hg1XI6YGvf0DhFXsQa0nKDPLCNsOELUVvao8UAc1u2L/XG5Fb3pQ6PIg5aMMGScP0wma+kZ+chVD
mZEfxnuY/fVcVLhuVrU7h86ABKKglMJGZNQBZNhrnHkw19mECO+cuMc7jin3LXoXZrWisT3mk/3f
nRRVHC6onEsWP4D1f3oC9aE78i69FRaoyvTnIohheXx2RVZO71twHOm1rbx+Q3cZZR/J/05OJNQB
6KnWW/lP5pUzlmyDgsE8aDJSF+mgxK4f8OjFgoZEAhPpggCsHbOnV+cZQlLfN9ANKkLwIWAdyhVk
tenMc5uVUYtSysOy0wJ2Hp7o5KLgBWEMVYX4R+khIMHDS3OCNOpKGbSeBoL9RWV1Bod8L9zIClWg
oiFwRBYkTZHrhcJPELGsGt3Dhsm3obvQzeYNP+8VwlHdptT32L16x7f2ZgYtlQG5F0GC/4hxHQ/j
c3Xx/ny89fBaHjBD0iRcBQ/0czhStuftqSCqjn/3TbMpSOg1BXtZvAd4wgCvXJJSHZ7HhwypSuhU
hwfQfL07Uk6xkQs5J9ILLAapMHRrIBSQzgtvZjVW7vB0daXARzIzaKfqSC+Cqg8THHp5sbYOoND5
O/qzZTTKtoZjY9P7+iHzI/d7L3IKNp8KwtuWiPShdnuxFhmIRXfzuyny9USoPRIT0km/UHXwgER9
KRlWNdN4k4EfecwGRJYWUMZQFO0Sx7ARZYOwd0uo2+R0oh4wtWSZ20qSV4msocZPFEfVNeAYsr5f
udjTZ7KZXtRgNFQE0HyDIbSudsrkss/IobZ4mfXEaz/nPlFGNqmktz8zPeXVRqek66wT9CooZCQe
RvQfgRxv2OabXT/O7OWXCW+10TZJKlIrTX+2NjxZWKWH3xejUQuK30vHWvz6q2tjMU0/pVEIE7ML
U0JIQ7XyeX2Z771HQt5tk0s4q2apbwbkNBHISeryJS8lS5rZVjh5YBttQAucTND3+zEXny79tUz7
SDg8/MznOUvxJ+1H5jUUZPIf0TlDWRWmML/pC9YEBOohVZA5RxWQF8jIwbRvU7BdHVsOFMFKLEZ8
Lcjf/vO5dxxQCOcMSyogXWNs70xS0If9L00AoVsqwh5QaXWfTEn/GscgVbxwOzxQzjGFz1/JPCJ0
cokn5DF5urc5NkcnC7Dd/ZzN3ZWl76q8L2luuCx5pXIa0klBjKR2/WRx+FzFp9JGgBmk6lJswHjv
dxmDZSyPe0g5sni7SWyAWgL701XCbEGReNmr6tfUumltHWFufpvWMLWcxV33XoRTWt5crGLt4scQ
5zt2SAMgvz1ac4f4f2d+3/+OT2yLt3aGX2Zmxcig7R0TBRYeSwFDmOpB9Sj4a7K8hxBEE43DQSRs
r96XNKjaP7+/IPxzM2LoMuy8t/sF9aCxtkcWqHGraJAnuGYW0gSUSrWun983xcIGmlRKpm6WIULg
H/slPEy+CSdMGErSXw6J9Yp0pN3/LklS9x74Te6gksXrJHWR+kEHKbk4xtHw0NgshMjvZZuzq/AL
Ap8o2AceoBSFR2mfv4cdZ9A+KQ+Gm8Vxnmd+0l1QP9VovfOzmS/DTxFCdf/xF6c6AnmsVG/cZr/A
pJLU9y8EV+3qqAwFlDIOnH3tLbNY7MzhMLSCVsDlsaIuar36ndlX77Rg8WjxZ/yxBUlsUqTI7T5C
9MSOthaldY5y2BZ9hz6agOxHVM26A0ds80juBSZSJj04jhN6V2zDWSeY5KbKNNsigK6OaBNgywUl
sYQd+B2v3YDZeXakqplrelQOd+Y5j31UZREn9mx1u3fTVEMJkeLhUA8ss2hwRVtD5QcxdaU0zrs5
6wryBhuT7bkjIVfbAI6JZh+I72w2r8QSZPTafgh4ko2czomWd/pwXQjrdN9ZVjf3jJ71PSNrdYao
PF40Fd3kHVdfGCL2iz8Yovzur/AHFN9ziHij2nUlpE5hpwTdfBbwc0jg8DXVoHInViOjt6uAeOjY
n6IWVOFx0irUQT38I4GR7JbBoWmAF4MEw5AJ+5u7KV/TlyEiTlyvFvngxLIVjackZ0Xx4Pego/YI
jmKk7RLt5VXhPnmJOziwfz8tAN80SKvaZ2qSKdGauY3yCFu3bVINWV8EU0XJslkoE6nOF98iOMNM
ym1pu56v+sLNt9omnwpmpGFolHq48kr6f07zgqYPpbwmR7kCp5yPIZbAqE+rk0Z2tTwlFfdKVlh7
vZkl9XNsDcIFr31Q+pHPw3gxIo3+cJ7LS25u9ns+CJqabgBqJkDLycxg/+6sRAz9PNx5zepZPWtM
sj98sQ87tc+Eiywi8QWNyNextYTay4auMThHk9XZeScvtYqeLnrlFIFFKZvJjtb34zs7M7DAYRkJ
s8+P4bFkCjhgso5Q0xss8vM6F7K8+2Xnx6M3FLG+zyOa6SPJbIgeVf0Yuny/+cdkEybsx4qCAsVv
lwoMsx0GFn2yEi4hQmlP7egZbdPHdccIj50iweZsmFaosnvAhvdCr4RHG7bKnDkwfG8jQYZXx4BX
7Ywgyhcxe7wiKNKt9oDNX1E1+IwTZoO8sD+fc8RwKYW3YdDi2KgwazTY0Z2GUS84jur1NxfvBeS4
OrzYvyAXErBz0ycYvqe9V9HXSYqmjUCgmfSWj43UdAWOozTRibMiUlCYF3X/NYMSJiUzsOgHpzDN
/Dujogidgjs19XjugZVf5gGEeCc4iQx+i7eza1BA25y0M6dpeT4mZ3V2CVo1XOE1yKdwG9FJUWrZ
snsgqhITaTNucbi+KHvvp1wC2nOQoHB0oR1rLl1tb0U4DhqRF8ogd11ZsTwIM/iv0dbIsHlOQqIX
n05IWU3r+YyOUHDLsakW/pCJQIOpToFqk8EenI4ZX89aaCMfv70gu48+vko5M9e6xFlYgzYMEWS4
qf6k4+Afvav/YgrV/lTzJ7lTwEjM/+p6IweIHy3O/TronZ096IbCIuNpAKX6aizqwzGEbRxgnKxX
32UQpl/y7Jk6Ya7SCKbdgg80M867txKXOmFiZI7vlwfiPq2wWMzZOo4mZ3JbWBto9Ts1uzW4ae3M
0LvxYCs1wLA2nRopqvLk/Wa1Ox78P5z8P7tCLopz5jJi+Xzp5+QV5d40Xnv9GIGAm5j3Wi1Q/HNv
0TWRQsGp4pgnIbGR3/VZ0QjPJhLX1V3D4b2StZjGkJb4RWKzCYn/pvsbgk5TMw8bkOV8FOJZedcE
Tvkz2DmIT3fcoWpS+h9SROgQFqpFHL0gpSctBFl9VO069a0AfauTOO8YE5KHveJngCSEjcBFF0PP
kCeo6R4SO1w7qH07JbNczCbBnsKnII9YPqjFSpQy2qtcUuh1zWzuX8u4E43p4bj7osL25lmFPBZX
dZR1yQv0jsaQXGcWKLLDk0qkwzh4j8e3tekBLXyyQrLn3RWKvwy7IwLpqWKVvFp8x6Y6Q6p64qOJ
XvVNGhysbrFtdNNe5bGaUh2oG79LIreK4pulYbaHYnqamqipz9zoA2aU44u4aN1kxM/usqkmipBL
9U0TeQ6fh6XTTb81fNY0CcH/4ej8vhhpb8+ms/y4LWK8TZvt1D9Drdl73813+9XZphMvuyIya0EH
io/rW3hBGjOzcnBq2U4IwfYsova2CkiRSWv0I6O70pmI3PRPE3ZHoWW1wbGT3Nj4IHgLxbzGH8sN
hGl/dkot4/0zWj2CYtNpl+f3gGVxHPeg81KFPH07d6UOqdvVw95NYJN2RjQ80tO18UREzYPef1qc
stVOc+Rd5NRtUzoZTgj6h7lkO///XxHwASDdgplqBCtW8i7Ub5kX/kP+pN2UOnADqyV4ml2Or7wA
UhH4e6+ApSaNCfJH0Rqg5a7Bccyml80BbaI0Ggv1v2rgkVnqCSCx1htDXGuEwpL1p3Ky8Nlb7m7L
DQHNScscSCeD1HIIL9kGS70WFvXjLUy9f72vMrhzCY1vaK0eHkh+sm3u2t/mALaHfgbzHqukr/iU
KJ7v3lodPasSfTW3OGkXbD0fK+4a6j70sKU8tVtJCccs9ctgpijuFdy6paWyMrssqOhNnE5+EOCD
q7wBxzcZOZBv/itn8Xyqdnz5wM3x3c8eH7wNT+8IRwNUvPFJzWhlHifN1HHTXxt/QY7PB0QBC5V+
nybdN4YLaMKp0w2RW1pAbU9s9TggFGEHvtYrUNB7i/mE8iLxfpzJMK3cb5rQISijWbymGZctenMn
rDOmoi7EaygI2VbKEih1Tgzr5Ykaj+/ZuhP46+Ym91sjKbxRMkXl0/HgLhQrZdNXzGRsqzshyQBH
/Nbm8wS3AshYGCurql1up6yiXlBPmAJ8Hm/pvE+NW0dHcs7mOyvuzlppkxkCbpwKYLiCPF8vGXSq
uphmeufw0T1/5TBxoBFgqYG5kB6sWLsk+YeItAwKcOnevOnC9R7dcHZVdbcPqAt3r0U84hzQMtRE
iuLEXEd/PJMMHZz57QIQPTLzaa66A1fevKk80uxV3Eqq1ISuEl3aAZpb+kXGenCrp3LjnMNvtVjs
6G4+pp1KoQaWtzLsu07DLLu84/xiTX4g9QtTFg2jGsUoz8orwGVhjBkEehwZ7P4dBRgNVC9BsbSv
qlkwRz+CkWgIo6tqLjHWhoVwFAd428NXB6mjCMrqpgnNyp2ENPwugp9TPvA1awisJMch+aXlD85K
OA/+lDqXAEODFb90W7ivB2DIIjMk3u07ZxhwxYZPu9biw9ICluIk5FrEmPS5zmR1IDNuAds06yVu
ZuASoUcNYumOLSMd4hnx97/I/YatdzfLCOjcsucratLCh0cG6SFm2e8DwXMdhg+4TFWBTFFT2prz
5jtKVofvSibO2aHNaSuCDokVNJOFr01aFu7+rbDV6GI7Yl5bXIRh7jokN8WSubyhYm2wlEVH4T+u
G4CCTkUjywcAONvMQ7Ij3oE60xE7DBa2nzm+v4CdjpHuCswGj6GVAWmmYqhrqg32H73ZIRzrmOr2
wA5yg0/J3W/iNFTKv3I617u9IvMv4UobhwAjGHMGgSzZGZzcaQn1ebqAKTpaqqrX7EbjRsaAbBj8
gvx611p0EGM9eF3bVDq0wdkRM7HdRHcBF5VWQpOfXhDsBLNsItbKAN/bdT2/OUj5HE+VVs6+YRVI
HskFcSoRj2DCYqBh+hMQsMBZ3MgGXka8gHCGYoTA9WA4WXKvfeXaYg9kQnCI8rBhup1EUzM6b+Ln
u+b0Ahup467yeiJBeKsS8cAiJpuZ1GFHu0OihGA8ea+tz7DSI4c6O+oRyBwV0HnULmaFc/hq4P1z
zNwjYmdC11k6MP0WRyRHTDfzeZXVrhOZFwCDijZarTy6/HF8rKKgpQtpEOWeSDyvo9URJOijJsUK
5dZwhTK1zYuJRrYDv5whJk+nON3MCgCkKEbpfGFRsXHb+mAWPiZaRTRteqmvC0GT1TPYQRzDOW14
PQq8ymKqJzMMUTqBeAkqpvKnm1JEb+zCxqJCo13wZFaWkBQCfka0FQeLEErR3VwyWW+arHHvM0/m
DVd+OavljWwG6AMlOY4y/NZbPpk3Dd3AAG4tLHcBLcHdOYiZpNESxcavcHiswOw270kKpNEtsyrX
NT7NtaqfOJeUDoU4qtas/wkASILls811CX8LuGSSJ1eESOjOLdjv9NEbtXWLhZIvIKFrcSvNsvZL
cFYWx5+3ZqHedLHqFk7AA9+yaiv0ya/cY1Yq0n8dSxtPVcn66zTtIJ+9s2v6iGiAFcsLaOumVzJ/
V6w5hCsMFSKlcGKxbbblZPWUHQFn328NPBBObYY3sH6jiMHgW8GgmWPKuH8BpQSCNsGVWmT4lCEP
hCdIlkJUndftmsCde9rGfG0ZaGjbexyzB3bCDWBym1nrpJO4QFBlhCT5sYU9TGvaPKltbDFGEJYj
7TGvj2C214fQ8zROJpt3prEb8Kqa6uvcd7Lig8MCeKFd9Po/EscsvXCfdNn/++w07tRjsrM3QvF7
oZxHfGrQX0WDnlN5ppd4+/ALUpfMwZOCq/0ZL67vXMZ3k/SbfOIOAgBozIbRp1C2iuNewg2i2NXF
2Vz2JpF7JAwH1Kvvwuho+VnnqNw6cQ36+KbuAYUEcvsg+Kp1GE9F0NTjBBJn999VAFvjdd/qr6RW
wk5Dy+sCoxUrEv7/HFyBMFln5izml2vVeWlwWQ7gdccQAmP6hJWYM8r+SybxCraGiyM1luH+kn2r
0ibjD7s+TTeEcoUc8vxEzbGNdXtRIcrbEQop7NGyqIi+Q6mA6CrcLLrWiLFCBoczpFeGwl3FxM3t
cQvPrzVVivVVx3bIb/TS0BhSUu5EWy0NzHS+Mo/0U4YNy3fQVv14QiDuYkjdk7wI1m/x9WVc0InS
e+/nevXVmgCSjFkOWfzIHvPIdPm0xnnIr8iIC80ukIYSX3usy4/6aW9RSfc9PSClgpIV96bMXGD+
f10nlpsImUZ3yoGXsO+CGntWd0TGkwFWskm3Ka8wozFHbPWJxfh/d2mROnUJf3owpvKKV7spIEUi
5yaApFILvJMLUkMGP97pNWv6HjAORAXErj3+l3wp81Vtjco/FKtknlKDF0ljXnllJ4ao0vS9xTy4
e1Xl1M/CQrslv35R3gKa3ezISJw83Wv9Q50DOuEN1F2cVwAsi4YAkMURgCZ0HteAHBwzT9BnTBG1
NCdl0mc5WqexmEfIJfyRKT9HvXs2MgluMFj7/OhiVXUng9gYoEQHbK6+WrJi5ob3iF/ylyoWT62G
S9OAM1SQONkbuamuvuvdjmwUM0nwJ7SybIWoW5HO+Bbfzj+6vCbWhL5pK8eV+KWnWfkRGGh0VqLY
uDQZfaeaYHvOR8dPPkfwOFoHUcQQIDbrA5EtT34i3Nu31knv2DjTDdGrxENKZBQhD/RNIbKysIQW
raWp3+fTJKcgBevKoeIVQ+wIJw93VjNMq2UrrczswUqmKKDs+1EkUPsk3UuoCmGV/lYvBHpqhHhz
i4kFP3YlUb14fQxlloizmwFqFq+90792e97yjSF9DnY4pBl1CstpyF6GRrOjG1f+bFIjzCF4ZqKd
8ggM/8hyWe2cibi6n4L981oym/ARud83x0Wym7ljAqX4QshcpglYjUU+15jmgwn/Z+KB9sMelGtB
N3D/8yPaejtFvlby0VYOEZIp2oAdyhOJrjotwoI7F0cGxu04ayZbz8OjHnXh23VG+M7mXFKrgEKc
cjcxZAAoWkq3ZXKj0US0LhI9wgtnLUzQsk0J8h9vg+x4NS63U/6G30WpPjrx2TGN6rf3AOwMJ7bG
YS6jrNiI5HDmsCD2D7QEr2How40NONygtZf6OwKlJALMWDJlSmnfgzlO3YtMYbEL22ypU0lRD7PF
Q7Lrxx/6iKXMvcXs7ZCkUBpjQxhU9Eb+y5Zur+SdhhjhV8wvIEe1zjTV1a9aJYghFls9CHQAhOja
EVlANROPDdh4Wpa3BMeERcZ5L29iuAPU3VEKcZESM8yS0infPloREpMjUUmQ+4dMNovqBCDTp2yS
rzhMzlET8A2r2+q1ctdXvdYb/su2vqM39OTCLD13wfnOS4qvbhMuPuh4scgakIk5KzChk5XEwWUs
kXPNAr2rKrB2vUft0tYLALIgrBkVgQZy4/mn6KrxIuVAIDgwuDH4dbiE792gM6FjuoZ0ShKpVAJ3
stSswXu6IIdU+5M/BzSRfwkPfr/USC5ES8v/BlaAOUi9UtDmCNNqJgl9e7rPmSgy4sYfDzW97wjU
w1UeImHSyy43M1+JudEI7OC7DuehL9DahHxIrvIAY94mRmFlfihufbbbY0O3qXzlHZBBL+/uUNyH
2EyOoSHocyYt0QIS1CeoVDbOcRh2QQtT2GWL57ri73UL4qUkf0sj1KsmrsCv5lte1GBqd+9285KW
gU2ANNE5g+mqq+jCii4yK2y5gDlP+SnPAl7q5KkhVN96tCbiJDDCm0XKk8yG33E/YtaoQikjSqex
bYwsxu+vgUbcGTsqgEpAlsT3KbDguZUfDvuNOn7vh6KPJcrFU1lTPUSvbQ47dTPVzRQwhX3AKOVA
B/WlgJu8r8PgbIiQ/dwFpzYZUJQubCyci1Izj465ksUjS82YtBnn3adHilNzylIx5wta5nha5pHY
QcwYsRGVs4mxkXLekwRzoidwtoZydrv1ikSfGmGPhwK4PMcO8R/xPKH6KRPxVkxgEoX6xPAFPt0r
hxtk9/N9JLaLS45QdrZiCcS4Fx4tER+a3LbgptpTSY7dmKVbceAh+lopfXWlctpfZGGEfzUDoTBO
XeI+axqsTqTErPp03lkM42PQr8YQAW2L6hRs6AsUmasY0dPgQFjaY8Q04tBZ1PwK82KLzQAnsz0A
22e40tTSIytbufnpM6WmeRd51G+rvIHRVEuobLRKBt4S5diut1VB8n4d2hwWmY0ONBlxFIgGnLhj
nyE42VqJPsCz03crstKvkvsrnBPNz9Rf6Y4qD3rPK8kQshFn+txiFsSX2MazHREPTcEU0/Yjx0Up
gP6JKElg+fNyRahEefvdRm2sHrJGKVGwmk688+bjlDcu8W3jnNIPRn2bhE30PgB6TJV91EmGY0bl
IVp18ugs8kkyG15VXxkOp6dOFFphedAID2VZZzraqDimgnHOZlIk8xbZ2bOq4i1XU9I+mdKAtAbB
NbKlXNZLDrjR4ygR0x3eq1FuxVIGf3OGHS8ZVqteoD60sO5SzcDmlLsvnKFiqDm1scmaujkt45hN
shiCUCfsQCqTtzDt+0afGrn3Ux/ftpuUtbnfNnvQP7/W/ssphIkv932zhyYOiGXafo49g506Kmci
Ldp1pxGTkhgO/Tl59eYTAEiDnuTIY+xDNMBjq0Y5QDXGXR6bHWoYE83SQHMlIGK4pU0T4bifxdib
weMmfQDbrIPgsDQA49x6ya7jMsrBIvZvNVaHQg9k3ZFmBTL9ZMtDfwQYHBQ1+eXb5wKdAav9I3Jf
KDDoGxMJJGL8cT1uDA9f72ZPewfk2KfNHszIySlQX3+saWj5XooQWfdN2urL4Y8CQCLgtkKw6v+C
SFES/vyLneL3c1cpMhkfp3/6Nt1cK9s1sTBZW9pydNfngHDGc2xMawu40VV1qvs1K7/Yb7cDyFU0
8rMZQvqHvg11vYFtDt4s+aSU0uQiNUuxP+AFE8BwQDcjLjxJVeOPd59MTXQHSoDibq2cWoWt+geV
vkyztUlIKr7GhBnDpDBSgtFbieAbmbMalHh91rfZwIhfwbuiNAaWSG8YfKVziZ45Nzh7G6ppwhi+
tT7K8TWTI0RqlCNYwfDRRTjCeBvVNO0VKCp/u9wD5puECCeQhTI6/bIx6W0UvaPh+q5DqMmQC59C
GNH+ThsRKO9cCMsrbY3RyPpmQdVyzFNUcLTKMy3VhIk3QsqanLVOeBHQR9WmxossZHHHY7acLBmU
LF0e7TtBWR0kErSy53ZWMpJykfXH5XR7ECLcC5nZbH9bRcYPCwi6HawKjUtfuagjEbJ9X25xQRnV
LX2ITyx+JSP7EmwssPsY61g07EgYtTqX9RX2CX5I2xeK1deNOcteXa19mhEEl1OvU+rla2A1opEp
La+WINsZENVYpmRI/ht4yAtfuSntITGRR05LFBIwRmKoUHbd1fTmjaMo2o1PrRpeSIixP0+mMZ/9
52aSNHvW6/JMydT5YHHYzZPObHALaUvHrKL0Xqdxz5hwfaNiQ/lWZ1hkqmrhT2VEZDvkoyKAemKu
d0OKBoiijQKkiHlNAoH1q2QiH1HW+bxz7I0tn8DwyEGqNe360AjNkks+Tk62mR8JOoUBz/k/qDFT
erUog/ttNFVkaOeCNVKwgswd+jJF27TBGOjS66SIALkDrRCoWuJJqxCgcgv0SxYok8hrm90/h1r1
8tFrd7iPH7y3agJV+59p+VZwRlGDyV4nS8CzyjsgvYK25byVZMss3Mn1RGsTCVAyJEbmO0vK5KTG
pJDcG/Qzdk+7R8Vrwf/co8pDfUjHMGZd7WTNuq7cMav8yKTBpdPx3JKsdnp4OSLZx6zTVwt6E17/
b8Lyshy5BTFT7Xaul3eTUW99cpjZWYOy1UtEvhqsrf7Lob6jiiRhEhiJAeiQf65GqEbMWxqm3bP4
OFuBWdurkFW8THmhYJd/mbGkh+us5tdUSlVU3tbZCtDKdKLRetlQV60Fw8fsAKorNkdrXkkmjm+o
dD82oYmoNnkNKZrIXWrx/vZpRvzb2va8v/waVeBDtnleORIc8R8SjUSJM3jnL8pnaOx1fNa3MZlA
Iu/GVXDE1t1jGZODWnEd2hDcewAEPB5FFinp2kx6/kPmARGO5hkF7DTOLZ+8H4AGgUzXKMGJuyqu
0w3h6JIkZHpzXLdIyOp6wYjPdskVsmYQnfFPU8HVUWMkojh6e8hKYQfC5hUdflyHrXJUg0Dyhg7g
uAFyZRaTP5W+yRKVaFF0uSsCy+K30j31qQigK6AqIKQ0TY4hy5YDbXRDYbGrzXBz+3WPgbPcda1X
j93LWlrLoB2jEiVDnAqXBRqjGNxskiZg4WNFnf42QYWn4YcGYRw0jUBKdD5jxKQiobn55pMXslao
b22EnzlJ6GzBLnc/pzNtVbM7UnzmLZNch2FeikrOB4q/kCgBT3sy/KUSd9jqoPYxRIBr/PTCDJ9I
KwztoV/bh83coQ1X61GwURZKQBAx8rMjZRD0jUgBaK+FP9oqQvqof/fdc35jiUcj1Bu9ateOB4a/
65Is4Jt8RBihz4n0sEFdDzfdrW0vjslO47Qp6rwxRjotlP7JbjhdOOrSl6N7LiiY9rVJ8kUlb3kY
CCwaMJjOzJd8yQYNi53HU23KdzSwQO1T+zka9o0hc51n35SEPRYPQtYK3ThUIb7KQHSJIAyon2/E
C0lK/PYqi4jLhy7+PurTeCtapVjzy4EAp4hcXaMr/tga8XiaLB13FmhRygfWOD4Jaxf9u0Muq2Gm
k6X82hpqUCe1/ysTURQd1sPoYVPam48D1uAMDoSYBGUqMAER/PJLPhJnpF4IgM6n8NV4Nc+3zfwY
qIa2dJMrOdYm0B0ay490PKvJMyU93sBx0XE2IUap9mvhUzN4xbMc3hy2SnJ5XdXTyHn0t1cWPA1M
yWq5LopRrvMJw/AxL2MBWFbhauM4oXX4MO95Y8dRDXwA5LVaTsQyIZd8SYqCmISYajW79Jzv4NWv
IgZtLUKTu/9I+DEFCnvQb00xZMvZ7+WM8A57wq3V6soBTHa74A88CefDBIcyVSlkoMSJr9MONIJ7
OcZo0ea1rlI9HP4avug+Se8Ur7+KEzkz3Sx4G7ScBcx7N5+25lWrc78BI+eY1Tw821yMobLq0X9v
pxo4B0eyHdPLPa6yRFZE3x6f8JYYaypbOzuIYC4OfO2GkBDuKEILbo0pX4nWLw56teHcaLgmD4BS
3Z4ndRjw4tJF/Gmr7E72DU3XrbnKltxfM+rxYs9fH2j9S6+qvC9rt+kaAyKgZSE6RsdSYZ/yuh71
B3K8rLBajwgRkgD5ae7/U6ubTunUEGbvSgZlvd0jU6M0/eCM/MUwyeIxbPuELn+18nvp6YCWOsZ4
cdQMkiGrM4yVUy0SlDPJHeATdAXYTkglYXZ4fA1BXvSAU9wUTun14BYa/kYawZWxno1/GxqIehFb
eNxGe6j29sqVZo6TCMz2Wfy5iULsHlsGj3fRQs06D6oOWRoSZFHzJ7JP6rRoiZ7a5s/5s21j4BUp
6WEs4wVazHSMcmQab3dgf4SzvGY5du8snmv2vuMXDPT108l6lTiWrMfAyxSuQRRzYub+230T1IS0
v2KNOfuoWUofBjnFtuWqOQQDqZNbG7W7WtyG7C9gw/aQ8wetY6TE1rgSEAwGbdfo5HRF+5tpbnOS
N3uToVT4c8rCyeS1UpNiN8yE117mAdaDJ9+61eHRIoMWK+y4kB0FrQvbsF92y+STvXQFlFrpbxvS
era1i9e0hUoPfl66LlEPxKDQUgUdLkD2qg53BSCLkU8nUaek+renEJ13gaR/7x7O4d/InaK3SIlz
scpwwobbZ9uUirteKRbkhkeZWMOKFea8rPu7TSRMA4zBRm8cbZC7LE3TXj5rb39TN4FoZr09Zrx5
3DdU18TA/32tJsfn97qhlZ9wEmr3lSiHY+qOcLwbcuSRrk1oKzgcwyDY9VppeYH3xysVe5iHJ9OZ
vetv46LiZuO+/ivFlQnVL5DQHjz+57fdHZ+LjSkqggoJ6hMQR05c0CtUf2PJ8+eZIxMW6YtR+wJr
W4XcrW91qb4Fow84W/yOazzfTi4vh7rxuQ97WvORCgl//xhbNNj1i1DEAG9ncFc7KTSTID4Z9pWV
pAAcpAxY2ZwOEpZxb2nx7PMJRYrPE5MJ7OIsGY1wOmTy59cNSKxox5nRYHEU9kOAgNfpimJ/zki8
z6m0wQBTXUYUIOiYhvlG5D0wXf/OoGTkgj6Dyk8WA9LnVH2vIzUzJdXyNZU0Bg1MKu5AGN7x37Zm
xcnFArvHVs/gPlwZR9ZTKsRLktmiFCo31HygIYp0N4Ipd+N6/e6tXRQs1TlShO2V3zmB1bfx+nDR
pz05hNAWmk/+WRrvbFIzB1k8/cGp9HRRkjeRHFTp7166RpjyXLdkrAzOW8u2fXQT+Tj9aUJFJAIp
nKkBgk2GLe05FhPOc3qoCFXMSExU77pVOUNCe2PYWqJE/YWYhmuQtpiCKMBFKq/Uw9GGzTbb/Fti
eEkwWNoMcAVj1ZZOpR/EP2JuMl1GwNNTa6WDB9xb9hg8OtwuZ2tpZPila+pReKbl0CiybuTVax2u
EbzGZJ1bDTCrbUwcai+u4c1FaqIfwD7S55aYLlK8EYPXreCyQhLsXc9njYpXs9xl/puWyo9lO6ws
5b3HWgd7ZnNjL3ZU+XFQc2kmTcJ/mxgFRw8hUIiOuK7saSKxoGHSr9RU7uTnnj9NDOVJJiFfpZHA
4EpFbbrzXMFdzfT1Cs5YLnWUPeTMQxt6xEcRmZp5YpdG8tyQnvoBnQR0p8EdIpRkM1xAG3Gyx2AZ
etS07DclKv5lDauTjWa2rQAdhmjQRW59l+PBHEoKBdD7oecAaxKxIRFRZXaqzVof9dyBNOJJW8wV
bKKQC7Cy6yzs0Fd3187kuCcap5ViceMEt6Ljo77oQe5xXLe4sphfCCxHg8vGOOWjJr5ltXGx0RqH
xRzYpU9YRcc3rUG3nmBAqsBGhkm2IaNDRMvpF20cOhVh0Gcv+A6/UQxnOhlheT1iHsbw8fCRxbFQ
j1xiSAyqfI46YigJltCu2hOODs6jaODX8Hdbk47BZPXmCpMkldiJLtmaI0CVE8Aexi/IepZo/zOx
ywpn4KGn1DaarOJSKYM7geD2eSKxMREqtFBWCBFvPCyXt2mbeWdteT0boGOfjfYPy3Bw355o/ehZ
OMZB5XFO+KKc7dIL5TwvBDFIbfn61YZuWCx4DQ9XyV68he6+DsRqqRjSqqhX44hcw0vplam1poxP
z69vaxDPnvZ6qTu62+qMRUevpJkUmXtNgXt+SEkTxQ5XmpgD9PSigaI/ctRd8Qkl6/MpNvoRkU9j
T5zSDGjWLXYWLVcX9I/Mpsmxq0iikiD8fqj5mVF1gtNu9M4dBWr1WlgA2j5RpRiAQj3LlCwDi60W
aO+24ZZOhe7ueM0aXxqzBRSOkDtlGss0YpPOY64DLj4+Ur3q6RCHsP8GLLWV+h6UKBLAXt7ucXrB
BS2vFPgv3LJZWFdAuBmMJbjyEgt6UfNEWK5k1/s6k0NF97MShe48MmKbZlBmfGMJIyAC09a5ii48
5Yj1tYsvKlH7QhDXlAcrxaO49Ge/pLwmp01ehuCxigzaanrtBWgg45eXu1kUwjwAxfaOYOvCOW75
mY5rq9VGrSCv3oDzOv/OdYdR7F2xkhUCEbvTHm2Cd6GqOxL/jGDpLReENGq/AnG3A+wxDQPzMyQp
JVgQCCd4aVl6b1lVQBfrwMU93P6n55S9Rek5wT18rikgtBrYkFj5JKNbgNTfQtcUsK9KNzR4vt35
cbev46OH8GnI7W/Dv6lbuiJvVvp3NHiK/mN8oqzKOwGbuWDD5JKoBuGCU4+5q1MePIEtzfsvuNTQ
SPy0/m1A1Xm8YuT0aQ5J77NgppaRoi3G0S8JVJtEV3MKae6BhlVnQGQePbAXsyxHap/R3J2rRPk2
MLGopSJWDQUAZsI7UxYyS5Ak9xT1CmnHNn766jEnZJPQ/sSYnVo060afgl9OoTAKQZELssR6upTc
UzI8c7Di6YJlXQPwPAjGcjNWauTi7dOFR349S2wa1LqYXVFCjv+Tgev+9dPiPTH6EdM4D2uTOJh+
GaBsiwxVvZaYbIu4Dk3CRgHPKErstQcp3ka+j08Ockmz/0GB+eKuu38IGzfUD09y1mkWVM9wTvKY
JXcj/SAbmP6cAPgGCQ2RtP/EVRh0/WBWrvxTPYZmpwGkw5l77eIfXcq3G+Zclcc+HJmZmh6DtKmc
cNf6fQROsz+7w3hOi2XGw5yytWNTZzl+BrBvrN7mophF4c0iWxqYC8J3YoqyEPAkAgXLwSdGxQCt
jtFRL7G2/tKmTqkmZHL6iRpFURAuNZMFzX2rDMPkA3OzZB0KK2npRggwwvAdFfSRyto465vbp1sr
wNgRgqAE5jCHIuCqmAnGbyhU53CVYGIh14qgYgsmh2Fm8GCWLeuGkWLa7BVVLqitvn4MrnSMEF8k
KeNks4W/8GdA22MDpWuKcWawPShAxteFGoMffHtD1EiQaLWov5hXRj6ekmPbEntV4GhZBnw1IpSe
9o6FG2wk7CHN6oUztfXpa1ycXSqFwqBnTibbncdmZm/LoU8FRSjWrpPoRPlYf9yuiEL87DxTDh2b
MeKKMpXpu7WCz1Nh0pZtVj77pBiRVUCBApqYaNzxWOV1HsorR0iwAjJXo1vP1z/TWhhGi8ML7PoM
RLQ7nmghBBbCzwc8YvQv+tiF9ejPaQFdVABk4Yqa6MK1/flYP2B4xVP/5bYGUMm6nMDQOqPz1dm/
9p3vjd/3/+HNtDuMAOqdWdgtfb65L5D79RKi0tIVX32X6noQ1tqxiuW7b+Pmkm962ekKM/vb8nAw
tVU/I9tH9WpMaRDBdaLP0teImIAbUqMyUf44/NQdHV3nzsktKHxkKwvlkkssDUsBtSrPOm5cW9Nf
w52bCZ/VUAxU5dbq0LU1iiRGoHMscgYvNIXylzGJiZfPWcsmUyqq9rJJ0dC18xqEuk2DrjcecIw8
RsSaOAVSzDoQCr7QzKh+BG5ke66y309cchwJE2n9+XDMg4uRuEMkNiGcc8vWdoCPbyjkojtnw5oc
GGrGz2BBi9IFCEYpGD6N8zkNL8G83+XWJxzvqIASnqvG2LqlhoI+Bwrx/yt5+XviCy/k8TOpWYuU
R0iBXBpEcrJyPBOzip5dtIdQgm5rHrrarmB/vvKnHWyMcSMp1jxfOZ1huVQs6imkRFuzyKou8PgE
jJ7MMGpH97TlcMkYrgGUM2f0f9VRIfwF+uweXT5EtP8BzAkJMaC13jRgFsKDXW/I8qnQr6hk6QxV
zQnc/M1kY2N2Ir6WzQQKIvHvBsJPVOrrZN/mCyp+2+Ca6ZpdP8GW5GoxYDT2XRH6+5ygAXbO4t3K
GhOWQEm8O1ICfOakpwP7T1d8imydmB2oGuwsbU3e6pWhq8C2o1+oUDRxYiPsthSdRe/ypT+jHFOp
RJ65NExeMp5+wdNsQS5SbzM/O9CWO0kHKlN749wJ3ckZOccxU3OzzuCHhDddcUzn9t2/YwY7e34B
nMVkpfdTPlgJhJ/vvU9rZQSlSDUcmUQT9yHxfW1kZcBSjP5HP8riPKlztw7UY5ZyQEVRlnQlnvF6
wzKe/WxXzZGuY7STPXd8ZFMiegkKzPKQDce7pO14/h6GzeAhqKHHVWDgobQYOyDpkbYvaqwCBI1b
UcJZmX7Sgvw6r7rEGBo5O+f+OwHI2AKGSN6HatQs08FgaM6qZI/XuCF8UCrvBijFyrQoy8hUQhvs
kxnUokOgEdgQfpY23OwQIHsUfbM/TMPzJn7v3SMSb15Zt/h0ggQqlkJJniKGSXaDEiM2/30jAClZ
7ZDqhSrQhclEjwR1k0bAbchCR0SeSdwLcgGoN/77opQj0KLTdjPG1Yw3xi2cywp4Af2nIjmDxZuQ
rmdrChRRVJ3tjUwcK9qGrKchumYU00Fsy8YggZFbctG6Dkv+lRfwNiwgZuPIZkYca8lsIn9zSOY3
2UFDjJiW6XkBZOoey6iOn1PyCpZqrfbP/N3dxPZKhNE9RgvJrCH3bqjAMtD7Hzjq+eHiFBkhLWCe
eQ9ASZ3BLpl2mdLoZLYco6lgQxdmiSPgjqNfpAnne8Y2KSbKc9Qtu7/WSGuvzz5rPOX6R1/KyaF8
SBs/snANEHBvaXTcdDSJ3uQP1oFPypg1aLoMILg1eay+Bm36LdUuwfmzCVCvq7H60NVymBbN/IQh
1I7W9bgnln8a1YZ/SKTvXZXt37QdGw7w8B7iS8I/rJceE5IyCGou+U2u+HlHu8ldtGS9h7NA60Rh
VzGqsgv/HYIhyRmHbl/Zsf6oezN8yJNGmChD7koduBMnqjwTm84NsOi54XoGsJcF+pTUpx5dQQad
IbjQXXZm0ssCtYXBsZ/aHPoQlsdwvNDvwELg4NWEJAw2VWpuMEunvVvN4Hox59xAoe5I5euN14qV
k4qgrNmZL1iLJY60eR0CElXmnKw9I2ryy+mVsCHxlUGgiD3F5ywACX64wmKQoVB9G7gxgtBjSLl+
upctC7SqdMALg2+7ctCneZfTIODs29sGURF6NRNNd16HbBmD+kgMrG5VpxgL3mHtzMwlA+mXZnKB
eKiavYcb0savOjMA+6Z2UZucxWApkc7uZ9bCWEgsDFRyea4LPTjlsglyPXFL3cCvSgI0F/emP/NH
oEd1MaJ40Ae+6VMcTA/aLrhVnBuk/vVlBjrlyCHDt1MXA0zcar4PxSGWUzT5x8oKYDF0LImKdT6j
P7hepKdVpRm+0Qt9oCNeVMDvl6Gmk/qHWUf7ScfjmpjxSmKoKmCD9Atkgm9+2GTdx89DfvpqLKyp
6cHuvrho+1xzTAV1csqgvz0Zls/Lr1cRsO57NdRNYFJPJOiHLXO48MYfaN+GJffQ03/caKKv19qw
WNihYXHwgDJLxSJLMSb/T77NnrwZ2Wl9ESo6+yCDJOAX0ZWodWj8NVytP81ImWGJixYbwHoG5xtI
FSq1gUnzDLfm9imGffIWilS/4dQEicDRdy23tCKin5Xa5iR0f1g0kQ9Xbj3NVne+cufVCTTEWXfa
SZhEIo9hdYR9dWVpaVoWTeUi8krCUVXKHjjWlRgkYds+hbGmXFH5xleLBSXeMNqVSC3XsJoQYkkP
V0vXwY/cLaN2qD2tQernaCiOxtO8bD+TNFy4jySrue06DpX/9g0NzYk/F4B/M9fTR7litSCj+bXe
DDB+UdBKlX/jdV4syU5YlDIYkkL07x9puLDtGejx2Ze/UX/shRi2ZHrEgE8MsimsypjZyj4N2TLF
JX4MsYecs4sZ2M2SxPr8dsh5FRXNui+6ijEp2hcVSVGhYPJ9m9Z1r75+MJmowdwfEhJ/GA8z3pNt
x2BGcRNEawR4GbodER9IG4zuODHu+g1kNVyLqWc4pbvDO5BiISGw7VBLm3Jql6TcgkwqUYgQ64Im
cyNybKcFMbqOzkXC0QEInnqWvq6r6LL8CvxXh6L8KnRRnfzfErMu49beyERUklfnzkBlhukvhOXo
1iw1dNiIU0lJgJiwFZIifPx5FBZarH30GHCXH1XXBme+jqOyQZ/0jbprkxacry6vxFK/rQxbD2On
J+LqZJsmzXbXELAy/dqtrNf7GtO3jnCkkFx01A3gm+p+n3USma2TcUn4GpvPoWozYMJgVVny0aRP
RtFH1NV3eWv/TNtZWW8KN0w7SsQ1NbdUxbHKsKOhhZcsyfSmB6USdYkAzjpmml8ooAHPhz5FmdQw
y+Zdxcg8wWgaOHFJs3zeqVwDDUuuiiWGsu6NkMcnu8yQyiMfvGXd7odNgQZHESlHgb7KMCmBow/o
ayzEqFVGb50StgDh7Ep9nK2LqxU+lRxcFtjFygHarXdgiOEns1hr30bLuQZ42wPmrTYO9/Ua511j
vzdgN/nD+SQ/vkQlm8vOzLL166DemTrakOr4spTZjRHILR8RyXJkqWz+ed4jVNKjGIjvlWYZdRjA
/j7YRSHHNCnHAf5HWwDz6U+YrT1ckKQktwL0+X5YIcm+y/y+O3qGZFGqWnaG+N81FrFyF0/G9Xsg
LcmmUBIbz9ii+C0mE+FO+ZTjIBS5UVEyY3MI6GRMV1waqvAZ9qjyH9T/rzMMnC3N2MQ04fbIVKMS
CGg27ZzDGMNDnxg8g0p86FPVFauIAqRVK3vo3jytJcjKdF5clQW2J1m/qelHOOp5T9yIp/gYxk/j
y6X3uRF7KD01d4gWAKgGKbVMEHK1jFqB/9Q91sQejb+uiIfMij5IYCrPKp2RQb74XoIAtd56g++r
EIwcSbzePz57CTBTDgPjjKWRIE+2ut4ver5E7HQ5Cjwo7J2dVCVkh7OJF0kt3jM2jdaAFNDYC81M
AEW+JmYgj1KjgpG9K4YwiGSLWkS4VDbpM4F0rgwsLsiQmpCEtbZzqdI1y7JtUDvpE1EakNVF6w0A
kZpaMTRDJXtf9DmJB8qmSsfsi8PxAuvXxb2dPQFCNp+YI+ZKoTz7GhudLVZ0sWZ6ILaInG5kYAz2
KEmzrWdBG9iArM9M3YsRCEUmhCmn9pJWEVvrPtWWDCCCJzjFN9hRiU4ZtDXAlR4IozBinz2/T24E
6RvShbB12JMGnEkhergESJIoesORA5l2rjbqw3lrL5N24sLiEk0tubhnfuiWGrT8TOY4GST0stWA
aWFwq8dh6auKt0sJrZvePxrkZz8lWdppW8RhwiE9rha8SuhnKxIXK6cxuHrYPLGm8+bd9GGhpbNc
2VCrnFZG+x9zujVozd9CVFPVjFb9m5q8igrPcoStZYJ3TM9Mi66cnFybrW6m+C7TMS+njSHSNUKZ
TEcmwd62Ju/qxfZ4YaM/py9yrrGre1vbRB4/HebyXAW5uixZPj6Goihy1WAZBRSoqoPmAH/0OYKH
88lZnh8o06UznbeeKdV1HKlIDJTJ9r1m3Gc9AJudoFudHuT1luCAJfRFxofVulU3aDxe5rnJaEUY
xWHdSR9rN7kyviVvcBkDimG/lzhErSTAUi/eCbFyUKlMTQQIvZ40acnPxdrOF/eAp7Ih/5hKsFH5
FO2d/QYj+iyCmiPj+G53fuLVKJkfdfHJUuJ3y90YvX0FU46Kxn1BOUOapZ/zMgMS1W5/zLh/Rpi4
pcWRvbSFPQMPUM1gauyi/kHzSJC6pNT7tiihA8FwJBnYB6HVtvqSOFieqST3HFN7WinRH5UImSRG
vgfo97AebwURtmhKxV7ypoddO900PLVzFgBJ53+NNmYHJp19j/LmToRZpeE6BRvmHDJj3J9IGnme
Q6tsWHZ6DSl7zdpY4T+cgX4OcOOLop/kpjd8GZSTPa4edvo6hQZ4keHJvXvivr+eIBILrvR34GPd
jB9vJYcIEW1GZ/9PYZ0jmoFhgwYxI7TC0DuyALPJnSBPbJfNZ5Klcrx129hQzJWlkyTOEe7VoJUN
uVqFEHNgBqCg9yKPgH+18jA3GJlTFOr4DP4ikr/jsJ6aHRw1EV5JFt4O7iRIBG/omCDsW3iUls3l
EqLA8p1EO556OoC3HllvKDRqnDOU5EQyAkUUUKBeufeCEwmf3o4O3RmWr3aNUUH4+WMZCk41Z6Uz
6xbs7xWwCeEaRmyazdtr3dlbKo71Ge+Z+e4Wwrs5CXlThKxDvGzX8bzmxB1ih8VPLeHiILQaJNcv
IYxA3mynB6B1EdJptZr9hAS/Xpf7iUWiiAhXWtS1m2WJ8Q/tSr02njU/EuYtaXVz0efwg3ao+uPG
R2TKR+wag38v5VaK+kHLqf+2S6HMsBjR9mu8C2r9Q7LrOaB4mZub0ozZVRPLNCxnE7S6Hu51eaaW
iF7zTkEZ5N5R2pDppT/Rh+hGcLLyipXNkUe2UvCotdfCBJHc+h90zKjoudDaTZjK0B1eYB78f1qH
4mFzdSet5N552HiqJQnhnrNlQWQO6lxLJHymi5ZeBSBpb+q+pE0sEFK1J6SVZ/+v7VZE5fzGH4F8
Wfm17K9qymzO7srX0e1fdMkXnMoFP55X5JxXJkBWjT9OaUc0RIRm72m8fnPQnBKeQ16hu2Uuj/iM
jq4LRoeoA8xDBiAulPjhI2Z6KXaMZ48pRF41iOCOHdvNicLj2lHwtb8UDWkMnJy0fDKwVQNhzddE
ZQpuvFlzEPjU5aSEQa20lUFGKg2galzu79PmDhpcOw+dqnv0zilgyFQrWsBonN1o+6ZLNriWLa4B
rTQ8kdcy4RDRJWLmsRwS1RrmbRa7j+qCYJsor9RR5h4k5nInu4EUgUa+QsTV8gpfikz+H0LNwIiq
lO8cYSrYGjX/bUinXNSJYKP43aL8LtProdZOMM1jqyGUvdQaKde5TiLMzjnPI7uw3I/eEnAnUYhO
0Ini06z4/QQFc4FPqXNnnmdJqIiQi97DI+5TfkvA+EpfHzHwPhLjtgasOsr/16zmFUxJ75TrTTFH
MZmJw/hZ0SCWrCGn7w7uwzxEkAhBEM0ZX0ose5OoKdNNdLUPcchTD8Tn2u5onwN4W5FmQIOMqqZ8
qcIQit2u/GbikVWqX5VtebCu6qsnT9zGXNZjN0hx0pLz8TYPA4KCaekdKksUmg0nqule8GfP+tMG
IYvGwp+PEmTtAVUzryMDIbrGcsjjwzwuzWxgmTmCPFs+UpQe5wwS0kxBNJeo5PG8Q46RSOu8g3Zp
cKy9e4Ea0OMUYMqqSrWqbprLOTCD/qad1yT8hYvk87p5vhd4/3sA7k4+J5fcX3FtObDfwbSDqI2P
Qb4Nwd5Zb+pXlkRD/hqfs3w+PVF6Q+lSz1wBkIRLwedvLwEu+8+upBcy0PPdhjdSMYZQ6gMmpngu
2UJNyJ0HQZiJewtN/5PwJIXv7jbfOAtG+w9LJ7zJsCe19re9a/ffF0c91t4Cg5xFDX59NAI8nEt+
WsKWeWdayabZJ9YVzG5JzTVnBpO6WoA15taM7smU9LJFZxijMHkSKJ2jRMGWCGI2B44Nl3RFGBHg
PeWD5bAYcTxXaswTtcOlIFXBGjhepZpXVbZJhUTLUXRyyyQVvvmDg6y2cU7q+gY1mQaqRPgqGU+r
7zn0v+caXBPav4NdCsGIs7UUyfticUjJJomDVf2OFFlOhdzR8oNaioF9IIHeOztqvhK14Xn6IlpU
uOMHywxNdWPbeVqgkfONx8Yx6qwaNs1TIc+2b/WZ8YhV6T4nfAwFKltwyjyE0i/TQrs1ngg2PmwJ
T9tsCkOQ5fDjxEghpYq4EKJgSRUq/NMM3LMtP2OwcOgAhFd5U+LQUqVveqFhErub7ovK4VQusyaF
rgddcHbAUs5Jfa1e6yTXA0Lmf6P/wl0OS+M+VfxKzPcamcjb2ITTtiX4/Bo92jidGj/2iIbA8iMt
dObxhRorsJCwd0IEJUHabBWkOnbBXzqWCP5IeKkIhBS4xMdnAwl/TUunBP/+mnj1bE/XqNf6zoHA
5ahCD53k3uCuCUdWA6qiEXa5LQeu2ZooQA9MamYttpyeSbSZt3EQEei8p3ZZ+sIDjwQrN7vYbA+K
GDcDME3IKvWMyuUBI1alViwWl0CluB1ihC60e4W4n4u7sfEYhqNHtZLe+PhHzXbA3c3gdIBdD9al
eielBl+KSEr09xAvpWWJeoke4y8z6UZIjA9vfd19tDOX/WGX7r9U0t9iRwfTIlcjrPXia8kRJCmo
7RFijkFoeyfwH4EFUaqbG6iBUMs7jXaIkXtk5SkiI5XVd95NOYLTMC6O9znUU3tTj0r6RUNFfoq4
fty3zswRkYOEFYU9w1CQEZZ36nSviz6Mh90TV+/RLMDQF8N1ItWKuM/mCY3At8rlSgnxA9uilkpF
88+e7JLRiGzAdeqnGY2ZmS0MyrQDBXhMOwQt+M4Y+A5qjKDHtYnHBomWCRW1h6UsmKUVBLusFGKP
zjvTpmmcAWmjIM7LYIldWBpGOIskpZiGUfWOXAMZgJgaUFkmRgGGXzJdnwrhH40x2Nozi8rypmnt
yqkT6M9Y/LxwgioK7bTJE3nYx5X0KeMrOCqHFW2peSvKZsusf9IC20xyXpIbe3CHth32Tfndc/8a
WccbwULzGOIFZqM9ekn6ycEnnuicFpXYbhTcE95Tk9k2zGnngRTuIKSsAXP/MFTZfsVl4yVizS5H
jssoHyQ+HOSKELHUWFaUhBRDKvhRYHh1Oh72IoYTSUftDuKHm7TGH8FenR05QsD55yxgfRMSVV53
QQmAwSQMegADC52BpKqIqMpqRsxH+EXR8Cc+b0EMj8QEwOTGQ82K8GtEq5FgQBTXYDo6jkF6ko4v
01nRtMySYH7TfA3pyYG7n2G7s+iY63+zos86OWU+oikh0TUZhzsA0V250fvUQJhnyrL01G1/BSpy
qTsturHOFV6SBc3xvjNgLcnBdG4aO5qcQ6HLjrkaoS1pQmcb4znB1V08rTefURl2DviwVCQOn2qd
KiX8Is08V+wlvtogyjTAJfTJbmgpbavov1TLYC1DfmbzumIaIhEMihJ79UxNxAEg6vm7T0rlHPmv
/0vbaoaCTacbhY70cdD/yJYlCjMBt63xg9NJycwGwi3msU80WTbtRyeQ/pnEvjYIPc5idALVI7TL
ao5cJU9K0dW+MNXkT7QA3RmYYB+aiyBGG2s0dUssDRq/NpbLxk+F4mjSzRd/vc6Bq/ePQVSQ0BW4
UUQ1F5kzhHwZAvf0uHWbAcyiWgf/n1+X1k7aFIMCRoozKYmVL2zIMGAAOzJMz8c5mRi5bgMyCZ+G
DEtRUg7jnOQ0lPHQBQ94LIfduiIKkCCUF3hudWmVNHjzh4LzZfHV8hw+tNEzwrCk0L0n389fe3L3
VkJfteWFSsdesXXkAUlKup3CHYikVDdn5f6EH1HqsQyNcC0thepBWj5kxIRZskvPrdS61pGeAx83
Jv85uBCd2VukzDRDEc8/oCsy/ebNbxjovBS9Wrmnj5c1QVPm2xGGJOpP8gCKGEnK8pkGm6n6ccoQ
tXWLSfsNk4LB8JqvXrCDDTUQBm0dpPf2xwZFCZTyv4IaLAK42iaTjniDahmitj06FNdAvCxeWYQC
iliXZYtDGSxMFk2xG/kLwjVxucJBkq/kEh3eRbh27hFKCBcI4joxSyHvwpFhSyriH7pUNYHKmupR
sbQhlkLaStX3g107OOqMSLKwINpMLvJcQW16pTh8mHi148n3rZCqQhmCZJsHc1ooOdhoKmFo2vjm
0a15cZtvqV8YbtJThWVvVJr+pnoaHwfMjCqxbAgRRTvch+SpPfEBv2dzZ3VM0mndIod4IcvOH/yC
IS6JJQkpcNXimzOGf+TLPIsCiioPpe9a7MPR8iloqQEIlA6izmrnTIA6KwVB4pas020KHyqgN3sO
E7GTRCZbKMietaJQBQXm/DU2pubwnLZmbzJR8Fv+rKkRTwb85vqKG6i7Q8+ip54c04ZKbYSo5urR
Q+29Eaqh/+bkXFnklGs+LylQYvyFQVfJo4sLezMnRcbHHVy1+0+IQMoO9kTFEzYZKwhXeFgCUe42
afPCs+HQ8z3nkNEvOUz7qynTlberZQSrpEeSKRPNXvy//OlxlkRrCpYdK06L5gT+Rlh7hHMEcsxK
CBrhdmLpcFIjFDegzSnMGGjMoL1KbYOVgPAKy+QAu+R4P3AR04XSSqWG8Z2WpHPGlQmMWWbqAhPS
m5g0v9qfATVK2HFF5BFolk58a0UD4De0XxkV+vePY0uSqhGAxjk7SBAV23q6w/hWGnS+4QYVnd3D
WLrOzHtIcIz2s8NFuYqNLLnOvIUeinuQWxYvXzpIm90W3cC+KtTj1WRYywK+jA6U0I+dg4+8cdsV
uGAc2tpHNa7LPol6OHaZLPYqN/QAMQpAL8V1IvIS9jUlhfsMrY+Ce1QlSZ4smuZt2kxlePn/RH7F
IZBwzn7si32cOpvbJkdCCLUlVFlFpee2kHEK/n20jKA9Lk9WXt47SnND6OWFbmicDuoJb1DBFIN8
BeExj9hH7/5vpT4Qn5aejhQm2b1Res6F4wMeguuqnq2ycJnZ9bnvZ/GFhSaPw1Ro7/4JRnw/iB+m
vcbI7Db68OWPYn+7bgRrP29pA+aEwaq6AfgMlZdpuigAEbCO/WTrx2uR7l5/cqBYJFET9oi1EVz3
JOv05TPTD7pt80r2AIhYPTWvWKkLfk7AeKJjK62iTavP/JkGboYOgQ677PJIZfulGbG6lI8h04lP
fukm+QQpE/EMb1ggR905YvqKRQoUs0Rz7n+b6xbmkGcCMcuIkWjMMDj9RU7XWhgYta/2XwX3Szma
pd5v3q6EBb9NPIXYyYxUeyaT3K8xbrxHBoXjBnD4zgVG+YRgiL/KLscm0u4+Zgwm1/LlmkAFwq/u
b3wCVx6cH7nmccp8gHKbAnUFRLLEGw5CQoEmPAdsHpMS+8MgTz4mymlR/2/JnNntp+GmQUOa8M2v
sfmDGnVSK5UTW+UNiYxGCiMQkwtRTU6HYcH0l/co46y4iPlnn7p6hC6Ojjh8yVFO09wJVjAQ5nOS
X80dd6gJCps2MvTnoKZt+qEW4AiK7Rvt15SYx3LP864KLEqZU+aXXlxTmyUb2GoJeyMnkNMcQ2j4
AEZyR+tli87lF1H4cu+k3zq4PBuOed3B9jlPQuUQD6QTt1thc9Jqnxc5OXgDB2sfnp2WgOqTcOW4
9U24tXgHYN/64XMd+vdSgjJaMaeYcZSlcI0Eg+RE625VqBKd36K4AZ+8aGEKHzV2LOKE5gvg+qK/
bk9OVI5AzSA8Hqm4ETYEj0TI+kLX5cJtey/VL4Ls6iuKJs5BxuHkmJMCxiO/9x7giK7dq44oJMS1
sCZglcDUVxtxkTrGHXYDRIPyzIa/K94neNAgaRXdhnfFa7s0BpqBoC++CzkmyXfG7p6R5+iVYmuJ
4ps4DTQc4RnA7am/FbaANGVH/YTjFQpBCkRtZJwiMi8SRb8F5nC2idB20tuIC9fh6/NeBgtLpLMP
IgFszotk7IlPqgK9VAUua3qGdHJCuKYhEtDhLL5wVkMmfHsA4HjTlLaubfGfhbI4SMi9M9Zx8czw
bkWRFTpfZx5ZpK1KhX18S/r1HDXrwAHgnXRJM718GLZJY/B93fEJ/TvZda0glLB37vaxvTycDpG1
Pv+kjrVnElk6hlTqL/9IjPSkKhm95Xz2hBj5d5cIGN/GTbhEBOspbMFE/2zn2iiRKGZ0T7X7F2et
rXMeX5rpHhAAxgFZokOX9J9TkJgbvmHlpYRwiQ24z5BneVm+FNg2XwvU5l5baBYywllQlMkuNwQU
h1uMKlVpvXCn7yWFzHJXRsgmok4Ruubj7hs4YXFL0aLLtKEJb2RdAKSyZkWwq5Fq9o/ZyiUjdeK6
slKAsF5MmATGlnZfmLa/armsepsedfUIY1vhB4FttRTHr0By2oyeLmZXF0kncJXvj/e4ng8oxrCH
U5BlxMpoguF1peDaBsNYZx3CAyVrIXC6YGPNP675P7EmGZTUSqozimskQ+0g2EBt2nc5VWvw9BNi
0cIGNTCFQLmNw7yuUZLfni14Ancs92WlK+sZQO5/25suZTD/9sc2ULF/mXSz7r3GtVODwhn9n3Es
quHDrSDEi+uvAxe6gc9MYnIloa7sb6k+9sGcmxA6fvu8zevq5ZfB1fzk27i/B02cLAdvM9LL/IrE
qhcUqZQwRd0yBYtkCZE1lYGZEHRLb/6/sap1SZ1R2NmDjNQTKyJnacGxAaaw/PRk/ISuL0jcouOF
lR/s5TwTg9vx6DFKV7cfPncgu68i96v2bC9HDFFSgUeHx6oH7HTQKPKfDcgvGXaKqvMD7NkVQrdm
Hf80SM2K2hNKj2eCJ6w20WNflXCjrGOh7cDNFFN7gLWkUJgRYuNKnflFETvj4t/FrFlQLBocDR7f
mPIcBTBaW6SCQFXRqA9XPz06U+8DB73eQuFWfWswLdJntRHr+H688MQDdytrNxe0HDAJF6s6z1zL
FhJNWh+Acr7D3qGp02Cng4dJS0fWdXC7x/ds3/jnEviQI9Gjzi8U4h/DwO3B7AJ043OrSXYhQhRL
1MBQyht5RxyQPQqzojcs6mF2q6NQ8yQ6ilkmawuA3/eW6p0Jjhr7KBkTywzvs1+c6PQNAaGhQRE0
UhhUzvC30gRD0dhR7I1FWMKdcMzx0eaQ0s/fifNLFI00bdaLgrjZ+U28zcIPIW7lH2WhjEoZ/caI
2O3HeM1DKw0RPemnwXoeXkinY8EjtQwZ5ILx/FDIlLBWi8ZLlELaTjQVjy9+AtEDF2ACOJu+DFSG
gZfD+2W2sHaYvICzEChnU6Mx5RB6vWRnRxIMBWViGNNXODdmvOnr7aMAMzpUZenOAR9GmcVVmeoV
Ktu/KBTeqmEBucLNy0JBXQu+6FXZ1Tom+7TX9eLouYllQ0jsRKgQdwrY+76DU3EFEgULrw5bzrPo
Bjt7xsLrxr648f2Yc9Ayofh2YnpjU9g+NF4Z5g/wGfhtfTh4V5cWjNn0WqqPH0Zbf2hixR/GgEWM
/VH2QaIZVoG8f2EN0+ApTrtG64NpWJMX2VnwwxW01UL5WRV1/+4tpFEbgGsMmZHitfrae5Zk015z
nkNOF497Ak0KqlRaH8Cl/jSjWdIWHWv2Qoj5O4tcgBze+xPrCXLUBD/9f0vQpLrZhJ3VjFcOKHOg
PykCOI37O4aeLYywAPnsLbbAoEx1wGhGDveCNaXl426aqggRcRIDKIpyLs/000jPXu2MkwTqlMon
VkmzJeR36/PFKlIx855TBQRqc1cYFHFlsP7i+F9oVL2Y5+UWXSGnv55YMd5Ue4mQ2W/TPQ3DhrsS
PRdGT/nbHVYj7XyfCHLx9vRn+9y/hz+H8lTizHMi/GzIsuGAlQi4CUF2wCv1IUSx6MXp1qXgE95D
vGZiQWmCGvBooTqGOxgA+IbSwT+MMSrGWmp27nrhR0ItL8cG1tE6blQwmwX7SKY47IgowpCXo6Sp
UgZVWYkDeFyyrUk4sjQdEa0x5fpM1P7DUrFCw06dtUOiqtN/jv02S1HayaiC+oOAJAy/qBwT0w+B
GMk+E3IhG95hOsKvaeqrtrjj56oSzqQqNE/GCBAahEr/b4hTgsk3dWibNtTVTq0Sqsn8ELVtpMb0
FyARQUwCU2B1bXMc8DEAK9Oiwdqh5Xyj5wik/p+kbbblgCaGP55jG1YWOIZf1MB6bWVFIQ5XPPyB
46LrbtZnFvkf7SUDo3NuZgLi64FekbVbW9YAVdCNWzQTEhVODlpDOzRkQiu5iJuyWGRv+RComm3u
J0/fcy0n9SdcSLe6qYGtJmeiJaPr14shE8n3MGIbFhbmw4uHAjJ3PKyFgRjGAiYse4Kx/soalZNQ
ma7s1QTgkuLy0kxCFUpVTVlmJypYJCp9q/5dYeNrUuIFHSc6VvNlkJ+1L2ojjp7VdYou4rYr+kGa
tkCkvxo3DCHlQDtSf4a9EJMtXyWekmqv3EIaPStw+beudTnbvelII8yk4ULGlynLBu3tLcnYg6Z6
PFB6SMHtuaG+g6zeFvwFCjL6ibcZVtKYYcVWpQEgUqYM4u2JLHfwuoOOp676f8SgJbML3ah8JOo4
7QgAjL/UiX42KQY4i3y3ILpw3QSeTHIPQmHRvPUJFRoeZwJbp25lDjSLFRd5/vR73Xi9PICcRUVq
IPeSrhhN8xMlgSJIvgui+kafmiKFyF0mtg/ehB3PwvJQV+c569vP504fMDX1kZ4gwEPq1aB1AXYr
1VBqvJNzM4t+ymBIgAryzyf0sWCiIL240Gms6cmdHd3LEyXsHxfk+uOtISbjxxY2/cccRKQhvLhU
48et5A7Boe528XcaolC2uhg9hcue4aTAHRl1Tm3RC2eWNNT17SJVS39nv1FUgIdKUg3w+AXKjWzb
IeXfH5ihEv/9RYpYx1JODIjs8HcCDQcY6BJZlZPT7+WT/luDLZvG7HD/CIYEB7FQIK0tPDphPlBF
hvwJyT9xGo4FftAUp7ga6WKT1D79QLppde6Ehgtai5AXR4C2L3drsxNk6sRZHtEE2Nm36hF3iNR3
aG9BY14HbB3hcOfdkuZHu++fMdTGH54IKv9aOwqDq9KrTChDOs79IYIzEk/c4H077Xs4gotvDf4H
mwLjCgZVyj8dEzI8dS1XisLZdbP9kzrZMs3PM11ttYNjC74M0uegnSBtbT1l3WZcPAdiDJFpmooQ
5LSU8k/bd0cZrYdiPtEjoH7mTML/gdH1FUqD/Ltxav5OGKeGmwmzlxG1XhWFWc5DA3cticB9ZDAO
QlT5RPpyLxeSl2WJ/lhHvOwoeHIx0eniFswxPGpjzqqTFpyFYvFSlb1PHesci21Q9MuMaseZfx5B
Hkiy8l++t/2khFY65t98/jR1y3mfYnBx0gqkP+jPp1/pQ7IRR3ZcUmWlfCssZGoilA42rVvnRf/8
hK2mEnonP7HFX72dMoZjsTQlspjkoyOOc4/ar1s8TkXhL4CC++BSSLhg1ANELFmIiCKu+E3Uix9U
HbNrYDLM6UenpGdmbtyvsh83zanQJmGSwJeXt+Z/alyDkrw7bJ8WqThZSbp/+JxXyaeh5jBIot9w
IBPgiDEpQgqmP14a67UD/lqM231igcvLqxWuCvxxUHNwGpyNBFtsfyhlPSDT5aNww4JRrhGh1pMn
67cfLRDSrmyvWW0qHJGE0tLe1MuWDfojew9coeCbXhWE6STKi8fxHxX/2PSdnfb4kwMuDnpMrZjE
m8fHG/yBXYxiGQFX8K7xCUQ+td6deeIlaDKi0cU299/OsKIbPiM5RQjz3JgzZTV2WauTeCOgs++y
NFZSd9ENlUr0pLNrms1ULN9ZL5XnrhLSJ57eocHN9OO05jM0h55cVEHjHeljA1/+lJ2VMdkJw50E
6n2mmRsDrHU7vrtmlyFoTYdzVCibCwV3EVVYNzlwba18EbFwwcWr8zXMTy+sOhhtfvBR3ud00rzM
BmJ4psnHcvf38D1ECJa51X/eOsVuWfuE0GGT7d+O+StgWrKBUIilcciP/1fz1ukFIFjcgBzDneBc
vME/MRC9/oAY6ziK8fMVlBB724uJPpsbQWo5UdFPM/OHz0WG1FbYtI9AT+JbH0fZCj40If4WG4AU
7eaMbbxVuh7tLLBEq9tPTI9Y+8KJXzSrH1naH0FkZDbIssgc2dr+VNlD0bgp0eQoLzVvNmrrmNFA
gFQwjm8NJ1cgSZZkkjsdsQJG+V05V0to6XBB2DorrB44toupTBNYa+R/kGnAMJ+i/1YY/MZ3wD45
p9zLsOkBGGSF7DHKWmBEijwQRpHmSipvG4wc6nOfdxRA001HcYT+iWnj+9NRQqK457RJgh9+xxpr
ZBnn/rkjPzAXLk3JEwA+tu7+R5Ay40hyHk4EdHfS83Xa/UbB6pqWNVN+zgynjgl8uE7LSM6KWWFH
7XLRuLzcIVNLLUYSCVkcYld/rWIZb6OSRvfA9Ptq52Bgl55TgnKkftUDzVwGQfMwY6vVYsJA51wX
PKJ58oVuf7U5bfmKt/8SGGfGIaHFVeYjW336cUbSCUriC5lwMlr+BJY46iHbkIN1zTzR+b2JNJuy
krlwQywBbSNsTdTgz64cTTsr5isWrVLSTwT6mFfbJPESBq5EVKD/Zay+/DM+p5ps9yboflgCUG6q
CS3Aj9ToVhgdlUfDpbUG3G77VaKvaqKkcoAnBTTrGww/s8KYAZ0vV1/hDlz7Iyu1tvw3PU8Pgzmc
ttBSaAoNwrYzvSIOW5bxgBBct1SlbrLc3P5ZgzGOYblXu6SD4KMoZ+qLh25E9UtDmd67uXKxDdtz
FS1AZct5dxp4ML5/yPTpZTBgj53qwuf158nUkrgh860myhx3ssN8LGGJe7FL8Vc1i5QzP48hs1kI
hXwUnVXIsS38QP0TMPkFlnFGr3CgGVn7pHioyryZvqPwdexcFKQkkW1c30YQnELU2zGz8OZz9FZq
V6I2r1H3YxOzdBbAbo+yNhfolb2G6E3xbeBhMkvFjC/S75Y6TjRhU/4dg+Yj32l1XnEAM/BBJuke
Xhl6cB7Imao2X20A/9RJu8ji6HiOdf+v9INrxNKQUXgoYfUASS7UQrXyNcy5Lkqo4vl0IzvqxtRz
W3XaT5enYmpFQldA0nwz4S2IQq3qE+MoSLH4Zz1vGEgVtDPnhCtMgYf4U0jkFhqG8yjrOHsfQRDY
tFZwHPyoLxD4ZgAwOzo9zyvfsRy0tE1sd4Oi8E6BNB6kc3k8YbM9CCNWmPlB0azAiG3jarYp6y3S
Si95sn4DA4yOv5ypMiW3w2wMKb7WB1qk2ZyeoILbk+l6D6UKjv2SR80TzuNO09udJ4QrWKbM04IE
/LSf8+LdYhPrqqJJ1GW+tzAv0mysHOJ8kD8IfNyoxnByvelZy184h0/tcPXw+sz4pyEbIkKqCIGA
qIQ0cJnRNGxvNepPMqER8D/1xvnqZ/IYsENvoFVDLRatKp2JDZt26I9dASbGAr2Gcu34YzZEi8CM
MQBPafzie4Ujt7ksWk77WybxMj26MhiVUYAiAWHYvelXKvsvFPDJgfiBrhZirYCBp3Eq6+0dfKRL
dU03PEr8x9yQBaZgZC3wpsJsbaLT/LasFNGlZBjPX4xhWRVU2wflFOw/B7hmC8GXkH48D54u/KW4
+TGaiVcfTKzpby0KIRSzkLaoAKYgYUO0SwjbdRbmIxhvnZvMRoXGB1OeRl/ivwUtDgt+8dUC4slN
bLrGOg6L08WTcTlZzMN1XL9FIlutSage0Z8oc78C26n7CaUU97BZN5IAImTVjuXk661/co337uqY
WiXzlPPDWMyLjLwd+MQwS4wVFaXNIqM5x2QJIa18pvEn6ze6Cb4q4jin1xJyZByB7Y2y5xpXHlm5
QJzRSyOpHTPvwOvX1Qu+abqBfoYW5Bhyf77br15aTlVI+rM6zDO5RaDb9VUxo7XgsjJQTaigFXvk
iU63OEze4vdy4e/Dvwj4/WqYIdUUy2UkGPBf/Atg81EmBWmpXqP5qPYHUWUwYeo26xGBO3ue0Q/g
Z4Dn5e3pYqmd07NegoalvsMy57M6vWcBEy9rossq3s2SMfV1VOGKDAmQnR5znJhW7UZ0Gsb/WW7f
o1b20ysuuq7eqVaSwvm3j09yCRr6Kct1anjDxDwipQD/ER5YAwrugUMkj3O+SX31Bo9h5/mbq8OD
ctYT3pNhIGgnE9kMVKmq2DTUWytd0Xqwb7Kj5XY+5jVorlbdzGmDRygALdpvlQYNXgIKvSMEwq2F
pqbD7wUIQcBPWsDGNHz4Kh6N05VIYcCwU0dOmha7FWH2zMMt1jXYeRh6yDdsdOGuEu5K+mFWZ0ap
KYSHbaUAD4s/8eQk/IqDmdr7F5KYzQGJwO+ZrF0D2LmBTXHlmVZ/lycLIyIYPz4hWUUwZv+EB78N
NXr5woHwqURuhan07v5qZL7GgOfpirk1A0i4u1XlJ0mYRb2XYquwTjch8tKXpuyq/NQ9vdLqzDyo
0z9KePJfetGJARbFUPlu/fitlIEFDP7CmMyC8Jl4lQ0pg5KqnkA/B5iSdoaJKAI2m677Cg+JmLAM
+JnjprrIndC6UJ29uDqR5QcdmEhkENgQ5BcGUkpYWpFPJ1wf3LUWdapLvsSZITCPhhftx4MTnEC8
7f9vJYiVsu9/yf2ODM4SBBZ5SswygtIK7R6YCU6MXIh+gCzf9GJZ7uiBC2liRds+yb42tTONaw7p
kzzGoMvpTERHKkhVU2pkSBSu1WNxwze89617hIoKsmjSgsxOaW70JntiIzJwRimWxXdYyHC2Q9Z0
6iH/+HEzuTN/N3Rz/+IddsHT9awsmLKQZLHZde+jpr5Nv4GwIDOc6rN0Et50IQo2gKVcBktKMfhN
HRsNaEJZ6+/iXrTX38N2ZQBUnHX3RvElWM6j92/1KEn4nMAUVgA/LvUtLEXF1WR9hEpbK4R9oX1F
BWDMIAKVrewB6bJi4q80iEPfYka08PL5T4QbxxFclrsqwyk6p92D0SnJRaaxVOi9iQIomkphz/pt
BH+BR7Zq8jW9gVBgMlIjkQrhqSwTrvDzpPvmdsWbFyGJzs8cE7AVKIB7wP8H061U1Y4/mRwQLTRF
sGD6SN+i8nvBenAbUjBtQu43zeRZluOK1WylksqdJMt6GmUU/6Nuha3I+rm555f668qHgRk00Lg/
B6jC8Cz72bn4SN+1LQaz7dzpArazS6ehsRN8dxA4Xz+Gd04u7PzdOb0hx/sVBWaLchqW+42GQYSr
15ln7HcGgwwbdjGAtHTkL3EFa91rZWDG/3HnpfzRMTw7ogarXHCKGImZUAxlwv+MUOBWg5ioFVAl
GbMg5jToPhit+BGIlQVwJZBSrPFwNvIffB21kDoKyBegn8vB09RO92i1f4um0ZkN/xoomOwY8XOz
EDH8G4bXdFRl6U3nN/fg3Ntu620p5+kV3XYTYP/Vx0G7ZQ4qQqpdQptqOMPhjvf5HtA/brwvi7lR
8jpl3U1wt3bSruTVcIYUi/G92MnBSR9D5/86Vtfh3b0AdTcL6wH5zOVfnLNy/4ID1+nujPxAEaXT
fFuQZiGBVRyDURh6rTX6YjaXSYuc2GEQW3MglT/PZ//2MXMOrk+jC7tnj6Kyj83fkQ2iBZaOzdvn
RbHYPgRlIOXCFkKa34HpgcA+HsxpG7cxrrHI3K4PO3LRebLRZowl2K/Aj3vALuRA+V900pJExBwc
2iBVOfCBbpG7jB6ru+0RJWwJcZHda9AqBUZM4Y86Ln7TvhHtXM/RFgPsPlKnpS9f8Zrx5bhSValQ
8c0SNUV2IwrHexqC+/aPVQ7ysoWzbh/WUOwULftX6AXx4zZs2Ndcl2rl5bjKfP8umDbbmoDOwKhh
IDBiwfl3aLS8ajwqAp2sXfKS8zQd1EBt594wjbqctMNHLhcv+d+Ptp/BU4omwfq+NXh5IbvP2rOf
j9/GDIlLAHMZ7093NREk2irF9fF2ACeiiJRdaLtfQgXHHleajbA04oAf1inpvv8dmgPVRgRsQeLB
KvQKexrOwGLTz3nSGOj+etRxxKQA1QNp6ZaZsVAN6DFGGb44VbXNA//IVO1UaJoNUL96YgchSh/Z
msapaV4V1QsK96wRG8C5D+FVXAUbuDx0Dnl64B61LRo7e8Pe5DiZoHBPzIvvERrge3J4C5L4oFVr
U+Uqsjiil1qLR5vw0WHYPbJY3xxPQE1HeziaQRdToU3KGg1MndYLoEIoASvxwjd+HSy21Yu5Zym/
GH5u0nqI1c7c5Lr2Pq+MyqJAUnmp+1xSEp6+FwUYomtay8pv8XgpM5LFL6bwpXDEceNdd1fgfMQm
JceuANUZXGft+MWs4Smfu8jjuEX60xZWtDBKwwh2HMKKKRBgKk3R+hyZb69bO/DrgmH6wNeBWN4z
uZAjbhPE6raH/I/BZukG+afI/sml8SVdgfV9Im3rCbass+lSpmvMToDoFfAenz9/PXvg97D4P6Hz
xlUeAOfuQSHjgreAT5mxVst/6VfEJ8LhZamvvbW6hIKdOIHH9saBPkN9k0BT5Ia1SJf/EyxeleJC
U8NeBeznWT71jNAV6TPWEL8AYfwgAjetz6nuFlknl+hbvIRRH/odfNw1PgLcFOd2mWkXjO8Zk4d1
hvXN1sorr6rM2QrytIrB6680VdmtKvDxVW0gHWkJ7n/eHmmv9NntY9VktDjzqtOtxUXlIZWMxh4w
D9P6ZKcMSZBCWZ2Fdfp5LdjWsnvHcKDPCRfqULTkM+cvtqzzGIhAQlSE2IAzBC6RvbqyDK7sBHLb
2YVHQEV9mxh19dZBZp6hxNY7MeuQvUzeyfarZ4i8OIj2yWW6yAyaWrjlPdMGtc1fO3xAsOc6675j
t+MYzVIp2MjyQebtfEwF407OnLl3gDJqRMgY5CKlEBgGfHiyduhO1fX8JdtUhE7YoV10VhZQBTYc
5Bw9v68eqmRBfNRoIjW75wlIoyH5VlFrlYS2wEkm5SAuZZUi/W2hUx1cTVri13Vy/9eeSGT1fOcN
mVg4SXW8CdPhciD33UKqQhhINiJh66OYX4YBuqBdVT1vSSZlKl4lilssyNSeFJEBpyARd6hR9rTC
U9F8gPRCU7LKG8TQN+ta7VfmaVWHAfrZFLXzGUevrgPhCxbIAB/y6ctAmxfID5Ssi2yhmPFb5QaY
nQ75SUnbN+cswrjE1dlNBlMo7VItQkM/R5xsL5j1DCUEUQLVCbBlhvl9sVWbxZ8UADEP7SOPWbrz
9scSGuHqJTy5VuySme0SqybD9hsB2tTBtZTxE4PfDC/Jmpb62dT1s3iH1iTFZZj27g/YyxqEfgw/
FVHARe+7uQwQdtbTt4B2u9ffrMAUR1DAtspANHN0/C3YZxLoPHZ+YdCFwrbBjHf6MgmBHXTqNUxF
UBfm5+gQZihkXzEPPN9TQqRppYHKn2phOsFbNkjg149cSqyEAIyovW9bqmPsNtCpnAmtHuuqRFzN
cYJyXAqEN+pTCJQouoDBCmi9vqKx2jLRYp1yarekcxgDiTBn73H6OpWtA5HneJOXUFnzoddzHPDd
ox74Vh5yeRUH+LIQnUR9yZbSJwOBsyYn02a0RdoktN2XBLS4Znz4mC8pKOiOpVp3LTqDKtYeq/4s
8aI/VCbnDzR75RFbpL5i2BFViVGEKUalLtUn8cSS/CvOOxXrVrtk9xnwaSKR0YVm1easfqc9XoW1
ZfUG3QJvRNor5+ync9yOZ/nxe8qXbHdTExe+o+cgnosaGANaMn4zxnw0tNCY0SVLT62kGoifarxW
4S6r1yyObhkg1aqCKuCh/XXiwRjPd+xeddQzWA1uifpnqr2g9HKdS/WPH+EfLC5pn4LltbZgr/p3
p4bGp8whCq8vJz2W3ka+EGf0mrG1648etGCWRlKS8PhTCCPW0YS3KZVRWH99lWvCCAtfOa8YOQbv
WC/BnmCRpBxICaAOfYi3HKZsdKlfp3NYbjs+ynzGqiLdPy6Z7GyXt0IzQxscJYBPwEGQ+kRfVKRv
gKqFfy1GqHBL/5Z6V6oXKu650J/5gy8sMIcUdE+BmHBrBPaxHYB2fKQadYgR1clhi43oQvhhnT58
BtjNRhg58/CForGje8OssarWlLMnYVPdjbnMeZGd5f3DFXEY87rbY4RIZrhm2djUbUYibFslYjnz
g9u9ZhW7psDtFLuuYK4pPv63kewavIfURravXLQnsWkRzWZXhqog/YbEqcs8LR/V5n7J6z/+yqUv
LXgClxIcO8h/fLLieNhSL15r76cukxH1slXJdky4ez24EnpI9tpGnk3CHVE+uLl8KDa8CtNmWhlN
VhdXnnPs2ppjQBZ+BFeIuyVXtOjKMS8/nr8uqoe6F60d670u8IXmTzUo5ukHr57S8CXKzjMUsoZQ
VKUQR2Eb1J5AxXKb0ne/l8TPw0Kw0ttowbD1vD/mNykicjyQqUS4HAAtpb42XJwBAPsTxv1VDDD0
54TVrBeNJzR3v+b+0iK/7l9Y+qipEZrbpOQ9QrDfAN5jg76Wltu6pMX2LrmPEceGNh2lEwtuU0yl
VDA5QvqZB/lFxbPgrjcTlb7+OEqoVyFlxcpXiQzjoZgctLVglqC2M0zscE+AqLM2LvRRvMVT1Iot
epPN/DPu3HvhuUsYbdJf3oBB0E7aDsbzUuGfFE7XC21Vd0+1CUfNEmh+iR/LZ+50HOako/Y9Ef9R
lCHPnV3MZjvyVdKYvU8Lbm0efgKjSOgsKkxhEktiy7KTFkaM9fnzdnvnn0Tsm3D6CUDJSBTTztGM
DmzomvYqRXzEAGFd8PAZ7JYpCaoDjOuhmfQTfsA/GJggwUFBGYZic/uYD2KHdO48YlPrNr+hz7Jn
bRCkqYm8SFoa6dzBZSqxHSZCQg/aO2vNErsW3wRxGOoxPfXwExlRUYRO4Jp1CaV7IyHG0FdX4flq
egUIJMwq0R6Cp6zvOWWgGbW4AxTrTDLELXD0waggac3KVE45TAqeMgBEseDQBByVzWn1tOcH1Rlw
khZeX0GlLH0Qiv58BgLhYzZQzVkta9xBMn0vTwXLP2kLOtDwI6JBCU/O60jlzZWQp4H1F5HZ3Ll8
a+G/kXb2o+GUNWZ+pmNDYlwsLu65bxsRz2AGaOJsnyy96NPN3hKRTtdc/wlgpwJbhhufBMXb8eYc
wEPnBS8gZUiI1pwkaFIFzudRIwwOrw997jFgFj0vngpez2QAYxfotfnX6a9XvDHjfAf10VHywF3q
hwZ/cUjYXVVsrPPe5hWl8WBDFoStgaUGm2B+FFHv0L7e9xSFXZyesvvUQ+2WZ+K6j/7nQYhdYW0x
YEUZSIoXhCw+TPpe+GH2O+DfHYArIz7w5faaxFKkOFtjtWVt1e+7XOS676JjOt7nLXd/beXwr1s5
yzGaUzWoujxfLETq7jLLzzYlOjmxOxw4gU3oFGiJXj696ncs4WBQ57Iy6rBK1GG9gMcJGXtzRCwB
k2h+hLDYFoOzOBDVm6bsHsY2izkupaCy+M+ge6uTgQiyoPaejgENWqWZANIp6gDK8AfZT8g=
`protect end_protected
