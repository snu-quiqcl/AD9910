`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p6lN73FZHRau4FVVDbU55VK5npWJ9A3l3NnyrVKkp9gRUsvTJrVEIDI5AGhcPVlJzqQ34dzBXFpx
wIKyyIg0CA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BUKmtqqTtx9zidF71+/yHZa3ECwGppp9LeuaKuDMoK0VR5mQDNuJXaVCAmN2w5n9dAmLlXyX0lnB
hGoIKUT+y3SSIqvIPqPCheTSMXYuiQ19pYW6TbzPDdVB9JnB7vh3NgLqyqa+g/2YAf06PNnoXS+V
SwfzHZBhLxfWRBtCdFU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SSR2s55Tzd6Ho1rxZyvcnfJWSZuItqujVg/Ap2/ljHzo96dSiyhBh4UV4vFcpNzNc5yyBasGN0vb
CTMWg9gZhRSLJKhzBqo8+AQK3ftX/GH/kig/b9fqHrdmgz56CgjHbWbeL8yd2jtGuYkGkG0sf/NJ
ocQeOhQ0dbCv2FZVWE5wpsf7Xfas4/w4OjjEHf6Sx0Qye7Xu7srwYt3P4syyEBgHrTZhvWu4xpzD
iw9rktc3Ddx/0EK+yRrBL/p8rvxhN1Gx0OiostZ7VgRmDDI0vKKe9R4/+Isb1n/6K/CbusvTmqTK
Y/j9hU9LY2BjUPOaOceuHCWmoB4IzmBVEPTe8g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Dwr8cPVfC/g5WUXU4QzkdTEeqGTXbRTHeTnZoCKUYhjDK9Wo//OEMFWAJg3GC2TdRHkEhi/ki2aN
0qSC7QDtNsjiorEz2eaGXgQ8myCJmQyBbyOTfu+03Tw45JKEOnRgoWxf0i3tejlLUotFCV2Euevx
dSLwnlTZa8O1F/M1ohbVQoru8rcL6yaeVaCqi26DLchfdNHq+l/t8ixM4LM3lh/EQL2BmVn1McUj
lhPRjpselY/vwqksQLmsOEisQhbUqHmgfwZBayfgCqjfr713CUYxddyw/mnkIBpVjLo8VulHo7qJ
heHvn/Md89VjZLFqMXrinpzpV7br+gK3y4OZ7w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lSj/MUZnadw1FeV6pQZgdWfaxYF0z9o09aAfY2RylqrTpJqY8wkncEsBeGqZE/vm8LFNBGTSwfhU
0jYASl6hml5cM0Kpe1wrbk8+wQYujTHAD642ml+hd/JI4CHeh+FIPf4uNeC5vvFjJgPtdrTtDgwl
5YTAlzM/n1RXVy7RMQouyRMB5RX91LA0+lr8zmlbASYR1Ecy/ZJ23G/Eq4aRf2Y1DX8IQCDhlA+3
NaDD2VbpWOJIuINpchvE71tnTS6PJXarg9GU6x2h5rxlpEaj3NDbAdOD4UMrDoPqHcFrKomHuD8Q
desEV2nbSKrXsjdkuKv2Z0ouaQAMQDJI3jGbmA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QLO8hCFNjwhTo3rtqaIQleebuiC8uv0t3YLeZPi2uK7/uFhPZfkk20Thvro6ouGpnUX/8E7gJZyd
DRaOxn3D1RSVxHpsHsKd6TvYEO+p6tZaJDlz3fc5+V/n0rWpRijLz8PFNVRH3BXu//E7zjiKnx1r
2bxonfHXZHGubFSHaNI=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ek7Lw8Qu6t8JykD1bpIfi9ibtmB5t6JrBSB030QOhViYDSlHMdQRPQEBNTQuot4Xm031OMpNmE/v
QgFZjYr2w1oFbcxibTmhWDLn6emdxlUjVO6b6XBHNhYTdl1h87GKBl0Y/kBHFRmJ7kevrwOYfxPP
SCNk95kUZlJChW7YSeQ4btgyJdbt7FdLQKuPqsU2hXZXD7/C+/30E4AadDqceDpjbt5vwudKDICe
PPXRLJhWW+TtUA7K+L9Smf0wvjPVoQBzfFH81ytsO2oHW53pfZ+t8NUbPVMYrCV5HYDoVtSbwjwy
ff0y302nEfx25mesbrTEG1rjsqMBKaQ+Dy2oWA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
eNsARdMJtVeTWx4qas2BZJuq+gDVP2w40dq8R2wrF1OSruHiEkVl9DVdqzqKUKdnyvlKarpZvybJ
lenQrVNxq6Vuh+L8zw8pn9LaMxL8YnUxa7r5SOhMv+tPkPSZY8snc7octBpqoL4VUuifsbb00bAb
j7kg9b2ZDVaQ+iRMaK0M3Cunt8qGkVqG/eeNiCrccfG9KMQCV23mQKh28PqB//qTH5if/AcUnh7Y
peVwmnXt6qkkrAOWKL5ZHL3O1Q4AxHpPskd2pwb3Fn3WOLyflwp/Hv7wiRQlbhqQIlxQA3fbh6we
5QLhGikuxCAAFLs3vPzAwNg64l/psiN5f7OM5cWjTD1XPVCjyI+9uWdoFdAZDkiWK8eMO7zrMkEp
fO4IAC1s0SBQXTeL5br4oKOpbM+wo/MSSDmceI+ynaGDJBZ5JhCpNVSjb5Xi68uOGwmhKgvO1Uui
ISvjtRTwFy3HMj/CRYn3Z0H3w/2ZkVaBBCA7pCqm7qPG9pH2jXb1rcJ/lV6cTc+cx0Jlf/4ubiE+
DIdObVosS37MW5A+SdRgJrvWL/79axQUkFGn0d6epORlGIbqm0+sH9xzQg7fr208/IRd94/mCSBK
8Hro/klAqvfN7SAOCXmMQTD6xIq2wjo9pz5n/tVguctup70SquYTg6eWPJGKbNqm8882n49UsDg9
bBDdC7Q5bBbXvwm1wQmd6exOlMEllAG/RUiC5T8yoJ/E+Kv5/OcjuY+3dy6hgv8CmSxvQHH63hG4
txG98OWVu40DS3QyzkJ1G/ayZNBvDdZrDlEcwSXjorjSwpnhBj3wf/G01zI5i0h+V+M4JYzdZ3JW
01z5l3sInSo2h5Y1oNaYiA8dEdRN+5ko8KRxqzsKHuKKOXWkEwp7sPfVFdsLNQQS+lCcj8wkGG8v
Z9wqwmM3JfpDf2/IXH2JW9FSiTCX1QUL7DyPC+TzN3lygdkgqZgSJPDPBy/GB4Vuys04VLRgMlaE
P1JNnav+SOExhX4ZYKMgKHj8/GNhpm1tQOT/JgOf4YzKrdMaqAvGZJFNJJIzFpltmS/ewpTQ1QFk
SFeJ4Op2aOI7MndsJG7EHmyzq+qqhFXO5Ln9ZSh/miomYTySGvwOSEHMMfnUw/RiwfeScx1pqa/w
nYSiPMdF0fbOYbHQCN8RBFSgOxuRBHYP+nFVNkpZRGoj/afSFpqLjLak0VswUvDXjYEUftylg36O
AAcsHwZX5H639A4ytVuOqDFadaFjmC59vL6YZ4IuwZ1YNT/ckpiC4rvY9a1wynM0f533uXLcVeh5
oyLMEmpZ/LCYbNzvp8wxLL3IAixVyQc1E5x2JLUGgDWkF2ePyH1YjIEZjqEtNOWvHfZTcGqaqbH2
nYbalkvXQW+uOV/Up/27/FffhXkqA6uqUwxYU/IKdTRnPc7WD4pIr/rx5sUySoQ8YzOrlQtgDwzb
FfdV/PkquP77cJKBgj6x76VOyH5MPpqW1lyUpR+i2PfYDB2cv4oBjC9SakxYmRuioL//SdugG6pY
AG6AiDh+hR5uVDEx/mQxfgGdCB8D1irULDL9uzjlq0OPKtbDwRXQg5GG4zRRkho1AmrKf/Cln0u4
BpB2kvZPLfxfSZvfSU0Nu8q6CYs5XtQ6YA96BpnRNOziVd4BsBG+EBs6wNi40fX7eulz+OskYg3t
spFqNfolvAaFuioNPX3FwermuXSLsaO5B481UzqZl35TxjLYN2R01IRCsXolFLvq+JD2hQGxBA5B
2kMk1sD2GE1wY+HvNfByg9MRVd+LPE7NvEP4PPU9/KNcMILbWMGwxziNcVZVAiPKIQArC/2SFQx0
RkU18Y1wckxrDhREhFZs1T6DzlXV1p8eouBUPBQxs027vU75zK3hBoAVqyKQDhoZxcEDt/w7rwBb
MrEEvntr7lI/U2os0TUcl/GxCL2QhIfRQ2YMz0UToa3kDSXRgGWyXduVzED/SL3NObTXlCk2SXXq
IHxbVS58o1GF4oivieztJoZvUU6lQagdbG9CqaUKh/3lS+hVFvfWEghri7wLMNt5nv4NekjKjf+s
uBfGpvluaif1VdEld9K9J6PNnTqAy86lAX1kxPDFflXgiVqr26y9u1716bq2mKbLiQUA9lFHK0pz
Y8UxyL8LQ4hcglEBv1vyngGpoQwfJQfaSGNIxtuMEfu1hCVXZsZRX0aDJsRq/NbMuz2aZdQ41QsF
QAQkxaooxOVftLFGtOq8JmEIBrMb6ZRykaI0S41EEU85Pd/qGmZkwuxbX8vAAkjUbx/0TIEtnb0D
TfrG1+NHORXznzoTWXM9tDkz5xTXOtvgtrysjTcVMn874DIwXYRpyvG1rjs6mQj76EevPdXmV5OM
lT2k+UNx58unOHN/jgIOGZKKIqVQBcEAPfjyjM1FhUXAxXsl8/i6yMkWSL3elPIWd/Q8qYE73GF7
fRqsV/lbpuy5bCFuwLjYbJ6ICoZf98dmY7C+zL7o6p9sIrQ6+XP/vzQ4KAaBQCE4dBOAqxZFv2qH
mErG95HEzOw06ikUjeEL1cnaq4j6+QAcCsdN8ytX1QrKFGqTGvbnf2uUw2oHb99CBF2EjDunkLWy
k+wfjyKWcVYN0IILWzERBiHmht8ZjUHJ6X2aFsWi+KDpsBhKFb6UdYyDag9K8Wxe1GwAanWGkj0S
cWhSeaHFXsFpi/IQZKsLK8TM6AAypdr3PF/66zkxnGGX36NTuqdY6i3zPXvW+/ScBrCaj7011fum
UqJL6LBMV4pahCybPZAWFyhp56Qz/Ddz/aieAbE44qFGXVDVIY6ihVQ27kIGKkGKa6eL+mybaULz
xfVT9riV/G69VrC6UyIfB3/eL78CbRRpzEfpiqGRXftiiAVFZlC/CTynzzKLdZJaC3LGeFm19+O2
wivNjPJsfAHFrN0PFQN1n4ppRTQOkVX9FZjtjNzatZViA8c3mcw2Pa6e5g51n+AsYgWvajTrVYT7
jAGKZMDgUiwWXbv8O1qV8ltts/igczOh47vzng/u85AvXtBsPb2+kPl6WwE25bQGhRW9L+aACded
uZnrMptS1Zj17jKR6et4ITCffzQ5H4EoW5riYH4PEiONm+5HRsFHUUXaq0Knu42iYMQcxXleLnsO
rizAY+bDli6/zMbJe0B/t2mnliMyym5XkL184UI+bTe+omist6WquFKjwyX8U5a/1f197x7XPR9f
b677guRqI/zzkDn9yYjgqGQCNdPsk2wzWrXnz37RW6pAOkpfe/C+OSYmzcgWWwFkXxuAh7LH38EZ
Q76eVr2Cqnv6zPxLysUN6LfJVedu9DB/2BqF9haIajk+uIdCHjzPajuyVck+HF/Lel9x9Z7JaLq7
OKDgmccbh5lkSPW4NFTBp8Cg7qSA3vMlsQV0wIh6JjfuP8cfWBbw3HcLkvqUsRGShmuCoDgPFTC+
MNWPA8qUCIEL3ZnM9t4t2xDZXFi2CxgEPMnKvf12sjudzFhbhgqqQhMMn74VCIOM/X4FQbmN/KbE
LQwXceqbuCE+kJjgS8nZUwIZQWObd32I21qbppsV8YGHAbi0jro6ceM4vYPQ/rXwgbpm1Q0bKP5B
OUbQaXTK7kHYEnzobpj1vxjR+oq6xUjHgYBY050U8fyX1S5KqqvJbOihd18Me9dA1DD3Bia1nypS
muvV5g+FpG35uxzSZbmIXQ7ffECGaQR5dePtwnpFAiy8R9buuNG+rHWGDBOge3xMA35qgOTtereb
WhThqCk8frqegYv+GDfEjqiEtZiIQ1z9qkYCy1QIhI0bFXXx5lzXIUDx6q/uq7aciY4GYhq0+J19
1mf2Sima8n0oKXBnjtl8LVp/upn9H6M8VFtoDkjhjnBiosWkCXt8ReBZYv+qJobfURxiKQslPDZM
EpRPzDFNtv63sGP6UPjDtsbco1wBE0sWs2XEuAhCpH8XCajtAlPRaG0eATDnJqSw4YLuv/ynY1eW
6Wq/0VlPFCA+RM1/QkGDWmVjc2p/xjdXINbjMpef7p2yHaKSL+g1ZIcmlCG0QskpNGHTo/jaP+F6
pixs9dttelF2UfOvxo/e2si3+FO7424jV9nuDWbIvSsROdhZ7btagK6dtMtUJbMoyIdFaYlgOAXn
6ypHmU1RXXrPG9CtEt+p5aeAQMXbANlIfGxgjupdmNs6ozp3Tv4tR9bGEK86wked5lN0eJLH1Zqi
kI5ofF0TVBiA3ekMirmFgQDYn6fDW8a8d4VhGKAI2NY1wEzqYt11a+oUJ/VrcRyzX4DBX9wuwmTh
QAdq8tt4vimcUMq8cwyn8o8Yv6+HthyUkK8Ni6PQ7yUsUgf2+1MEngmoAaX3xxJVqhNT6Is1sone
EPBIsPVUPT+R9XnGFZHxau1jhnaO/6mRoSQxaOUR2WTLTDj5XUt1pjVwIg6rQ7uVVz/ey1m0LtNE
Itxu232MzMArwKztTll/naHzOvojUjFA5t18ZMOYZbjYo/yTuEo6djKaTxD8A8uWK68TiSmjR/hL
c7HlFsU9p/r3sUW9tfSkok0Ay5aGPzrhkIoUu3kJUHgrb7ea9TCXYBHFJhlP03jkKpVaNgrWfm5g
kppoPYdOuKOKd3fjM1q8W4GD1uMpV60je1vjQ5cEyENISAfi2P1bX1W6j9MvUJEtTJrjlFl/DaRs
1qFMApOu5+9R6FDAPcCzFJLnHEWl2+9r3k+nz+ITQ7B7vm0w7ScYWdEMGqGpQrVhs6rP73XMJ3ZV
c2DMOX/ZYfbuism1AGiKPs3aqq+7LmVirYEHwGT+MZBaOc3hQaUFkU79f6JNgek7YKzANd5Z2E/3
KMIWcxe+ugXUbB+B0b+G4COjd8LDwctN77H4b14zw7tOkh9EjIp7aRpWmJT/clsfJ445uqjHCR3P
wk8c/cOz9hwwijb2B1t2wHVQlFbbHjLgHFTznbuzgk9u7ulcU9EI5gRyTs2+8tpI9eVqMwtuJTL1
ZuOvmUySLAt/8iuM7qelmNJUXWGMP/F/gq47DMpUwpMz7MEqury5QNaO3lDf1SyUMcL8UDJXxMzw
Jp4WGU4NRnlCOkTPWQ8TS3cZUYKo0T1VT0kiNQJT0HRXILpmAEcsJxWLVn8PKceXgG0Apc224QtF
p+L7LlF4+QmIBj2pnj94vpCLuYoXl+dymdiXiKGPMZTl30potaEBZ2eZltfW0ygYXvrHCyjAQN7f
9OHdse8g6SHg0n1BmWr5rzLQ+aF87Y/taq93dC/f91MJ7kiI9d2HNzhYSBgwidZE4fLXsCFs/GaS
cRoPKTvTZpROjYidqp2hcOMhvBRCR/eF/DMqGb/SMRnjeqSQZoPwR6qTGlC5wh/Dy2JqJWG+X4BN
Efl8J478J2kPxQDYZi41bsag5eM2iyuZAKgTrpqL+9CNDyyHoRkLkyMSBvrQDswq4fn6ECPWKr43
TMk3DvG4jiAgk3hkx8uWYi+RUOksS4Ez2dxWmqetcxfdcEp66nRtogFXfUkQSe+1DGggEhHEn/UK
3v2r1Ms3c3Di1v8V6WGWPCMGMhFy2Lrr9otmcDm2r4rUkZVeR2Qa7TzoN2lmUjAXATWOFwgMexTN
D5mSA6WSdaxJyF2ZMg+7F/jxhx9xO+OjmWJ+U/r85iqCbrWieOONOrwsytr3Psodw67HTdporhzx
fxGySpQDvVZVMOARCqBQ6FH5fDtca5LhY9RyW8Ih0eIcdh75peW2tTvrfwEY5RA1+rYPicXdkwqi
cUFi9aAsi/omkVcnV1sjza74gsX13IXdovkKrPzZyT07rCJZKX/lY8v78GG9kf4OlJSIVR2kk0Wo
C0jtdXCEKBDB6dlm31BDTLE2wgRdgFN30bwUNv6a/kBEb+EEfB2y12xNO3UsaaRQIXN2DlWKZ8ML
qALHOvb1Mp0FbNij56zUeD9aaRYPqUupujVA8B2eVxS2TvkCdCDmY67tYWjJo9P42u1lgDxdttzc
5b3tqgS0wURerVZwrfAtHx/m05Est2mv/yysO/Suw+gBZ5tQzUTM4iMk9npWonIeKGciKWNCsHQ4
wPdAlX+MOZdBXx78MnNLFRq1Hz21JaNECB2Fy3utvOCedIQsihjAAHnN+RYczxZ20Lmf0z6/ewqP
ETXDQtWs6Rg1w3tpAP6ZFss5pgtQ/XiYtxX8n+9wgIKFQOEs4h1wMmos5JYgk4mEzUCkuu5r6kzu
uj/6k27xpz8H40SKsl9pnX5ZKDsWG8eYTIm4cL0WMqwRNFVz3NJJGHYQjENzqQw1YiQmTYnnX/yX
keC+Gy2unfEL16h/EKFZbrYQAnmy5h6ZO1L+xQHLboX31NdMJOrT85GvIk9WHeyTwLdfEi3xLb6j
o+iiTutHcNSJn00mpJs037T5guccEjo4q8fnhJrzcVRoKHddhGbiquaMk6sKRIuWmJb05Pv1mtcU
U2Z94xMdVW+P7elDSRy/cndZnYzlqLFlOMoKhWp/q8YBuj1ZRM5HzURDZvuCm9GqJyqfzHMFUrvp
rsn8YVyb3PWQkhdcsSufx8F36GneG4Cz66aMdneyZpA02SecnN7HBy0N11rXAd1o51dvkQTSO9Z7
zOp25Pq4pMF6TlQXzBElXNFznJ+wpUWe35G1i+kU1UORqsMTUTxiCYSxeuph8d6+Sw/E+gKt53Kz
OhoGmE0hj808PMJrnVmAQVkejO+2vBxobGZ56LVBxYRMzQxiu3gUnSTtJiv75JZqDrZanujfHnSh
pvvJpd+GQVNw+dCBkAubTnSS66luXv/YcYAVru4st7LHD+Xa0Ion+KFbYfbbk/8Z+v9zk9Cji7GK
9v1NAyDBph57F0z9l3DH9GYrXcwK6957oYl7ei8W6wHaMcf9s97zjXkChK9Xt+zZZkmEuzUvM99J
J2YOAFTAZZNTDWXITt1XHH8TxsQDRy2dlPfyd95tEV+IFsAMKOD9GIqwEVCxC1PDdDRTy/JiUquF
NExcyybppUSBprhzhX//AAeZ/DJfJ+UXcsrw9VLynwnhFdVrGOxEjSs6YWwRJtfbLajoVC/xdC5b
qh+F+/go9RY7cGPReAJGyKRetyrSvlVj1xF8etwhMs0WJkA72ozk9I36eq3O0Vg9mNyCBxQVsmuz
j9OYeLau2EHfChBkzpmbthmHSve/fMhArmeqiCZ8gyi0Js7ejbsBhPsWdioAWTjdoltf1WEOl7Th
PUBu16rqoHJQaRisl8P73PIRT4YhbrY4s5HfW0NabBX982yhTlrX9otX+RKZekknoXGp8JNaTn6f
xrLiLZhwAdAauiS13qCLt8yTUDoVSDYLYiMc+sUAxD2WnkSNPN3kiUSeMdH5/KVCRXPttDixcjlf
aN41jaAtvZA6SfTw2CBJLHOZDuNcLlCGgY/hgfGhsRMlunf9PMbeLd/WFZIaaUoeTBmwRdzN2bGB
rlT4CJlbtL5NdF2SNrwpiMegcnjC+P0wJ/NvaWiekB5uUv7/IrlQsZWW2TFT6nBosjvdZEUDf8eh
do4OOJk0jVZS9XSFAbEc8GsYafpxQZa2kz+WPYkjIF7mf0DnBSyXrSoXK+cPvWOn5OnHGzvibsss
m29lXf/xe6egAShBd1tG5+wiK1HyRvYQZ5LGMWv76HVW+0TfomEliJixj9uLzhGgdn+gLipti/1W
PxF7DP+QfMdle98Pb/4CuOSuNiGXbkKcZqVyGDHwijTLlCQCwyTqKSRIc41GUwLiS0JNkUOdVxKW
FniMK3tflC/TnA6qfYhu+y2yZPsTzOGqBuH6zHT+9uX2jNu0SoHsJ1kdJmKVISJcQbCzaMU3I/G1
xuiKSa/TXCPTbX8MGh4Ybyq7QVV1s8PAmScmdiU7VyFGbNBA2M6l5Ao2E2mgqP5hYww4Vx/VzMnt
+GBTj3JtVepZU/QowsHoeEh1uRN4BrxBcbQNYXVgFsFiN+9kRL5AZov7HlFCQrDCtf6GFv/91pxA
giBpaer1+5GTRubm8rO7giG2WcJu31DhJ6G1X4oFArquWiej3D8OmSe3z2ibUptI0yXtdirzsDGW
e925xgZ/d8AMHBmwWhCAQS6V1wfzUNX43dCSBXBUfLZOeruSqBGcbzNsm2qeuoE/3WVcHP29r2oY
E4pC6e9J4jAqqb0sHDLEGfCWHPPc87SLMbgZMQiBSLmXh+sh/9REDrGR+VsLHcomKG1XwXd8n35N
3UeCwjfKIhCb4jHM9q9XnHzOmXvQ0JsXgc7XQswCUzrIf24zATLf0eo+lQCdf7peI9M2kFHu1slX
yDP/48bbAQLlXvMWQl6eLHVwno2YRl9pJazWU7LrC79TLQYylM3+BoQO+f8zjfpniBsRPamR/jaw
CG9gFGKJYkQ9rsVTMhXLDkxJsK3Rlnb68euxB9FiKuNr6Mioc3hAJmy45lqJyDfal65ZllnHsRJm
y3+VroLAEXCN9tGd7HMTMHGDTrZ92+svWWsq/V7yMlzoMkjv7SVJ8HRhY6solxl5mmbHoBXoEGU+
XJiVD+4T1BfA4SszMXWol0eCL4mrQ6CsryxejGITmH99VqOBS8ZwirREOH/q7KWOZR6DlXRq74jY
1hdHYcg4R1qvhXALV95yG50Z5YBNfMS7MWdWFkhK7EbxDtbJKjk62aMBrYxDnz9RBQkBw0GEHQK6
sq/Rp1ShxA4DRl2MCmuuZOhYGSymvDCRqXF1wptS4okaloJS6lK66tkeCHPX14+mNFKOMNssSFra
oTYHjRdMoL/HeU2U3LWVjihzzOPyIRgHDSF+EVzIIayX1edl/r+U27hwUhY0PXSm6pY8vINLl45e
V4Kt3NRxopxJSp4ai0qjrsm9beL269jR3qZ4KzuMMbX/FBG4oZuEdgdJS4rQNkJy1mhQR4hYa/Mg
Z7z5w9hjE/PieBryCRis/NUwsXGj+3zW9/u6vr1FCLpyLNa76vwEdNhiqbB4PUgtnu/TrTWkcQvP
W++ddhTtzbtYUXcyWo3Mfw3MD/0jitFKich41igu0ViNWKrD80KcdHahfv+KAVfFOR9vU/+kMsmv
+FmFOE+t5HCmf7ogKfwHJN4boaN8tKg+ESOp0MtHpdWGybHwyIQRrw+bhZ1/LQiGAZGPmu65TFxA
azPBvoNs9e5D3Nl66poBdGcMLobWHH1ZtDfA12Bp7l5RPjFcsG0x4AtnbWDhl5e1MuGSdMBwtaaD
pL26gfads88dzOI2oNtXhWDaHHP9CsuGhU6Xxl6Z9QORQr9Cnbr3cgAXMjqew5vmpsTz1XxyKjD1
bVJTHs+SSIN1WgyVu0rvXGwH+++r6M99BwrvVY+SxkhgLxktChtSGlZbOAjVvYF2J8lDd5aRXlwV
5kN6/tPaMBRxNNtt/2CWulHRlrP5tf/dSVWq/Bm+7jmu521V7mgjmHgQaLCk/mfDrveEYDTClBlz
gPqPFnPK77G2q25pZBhUfuuGhB+3HKKvPdw6JtxZx8tH8nvHa6ySSRDcwzO2EYujGk1kqXuq4cVa
FMD3YEVYTH1gWS58948CFm+H5fFU7hi7gdNv+Dg8K7AJT4VHTiZqiiKohos8/2Zi67MQNpFWXLQw
I+koBWhz7ff7wtzkUREmzcWpmLXpfIALRv09hUPE+vzsOxKVn0nqq8Mi6Z0yl6FOYAo5D1CY1XMH
KKs3H1sIx5FAImWHuSkxyQFydHqXxrYlYaXPlmDA1saw7l0y9vR5hd2wWyT7fFQOn9706aYZrx1E
ZeB7TYWEjC1H0Hi9dDcID+SITOeh/0X5yG/aFwXqq+QT2573bNkk+P84ov8w4YL9nwNr1evIWVDu
a1/qZqTQIt9MbMd3sn7cOHbmOX0L4TCUauxxQp+IbjnkEEqBOhijkRmzno9p3eAQTezUs6BQ4WXD
rElJ0lnh2gODvhGk8xhlHchqVfz5LyE/+KrDkVLphyzjBLSFlAkK2CVmvU4fnKE1QhKCGzSJHPRz
qMqoE1ppHYNg2AQdNPLCreKthxuK4cb9QoktYO45yokVKh+4Fr8AUM+zChztb+17GQFDFLI6zLe8
SGKweQ+4HD3QoaTlQDHpsvsGDFimUO3WmBNAlwY5zGm5fk8kHdd4WXLclTG4sDaKhoc4IccrmACx
OiQwkCB8PylQ8XR3rAAPozX4yPZcOtCVt5r68GJ4TLLRujPPkqrS5vsLQtBNSKCdoIbeTYvh3hki
SDH1iDrg16RQOPpQmxQPBf+N1GiN1lWwWcHCaGfBVBalIhpFkeDR8accUkyWMAbLBizP4ZTgOtFc
y2xFdiM8wz2b/VaLCT+WXGQK+g+zr5mnKVlsFQ1FcUa1SCNGsnj3rqgubylr68cTW/GFG3DUO6UI
MXCaUashLKuKU1R6wo3T6JGc+PraiG0zXt0pumQMGI36N5XeO2JYK+klvH4McB48zKrb4gaG+mln
lBhLi+puTRsSyccmtGxVCHzv4/8tfuuJAdMpQsJy4ys/p6etxhvq2VNpGoz3ste54wCXzZHhPl1N
w/LbWa9XaFYa1hn1IzIlYvGafIPsGG6svtRi5kWK+iK+VSa6CEdfpsU1PKug3AYdzJbvljj7nmYn
O/grzdZoAqWRruqrxwkQmExV+fujauU9Oba51pySXq8GNY/DLvCrhp3BJJflIwY7w2N9SPUoSgqT
P5Oe8uciTFfuv3XJdnsO+QpzdhrkeXNCDg7JN8evYJXwyUJ1Z0ale3PDK9Y+yKNKcZaVWFW5woT3
ee+ZvXt2+W9Ywfn8A1j0kBvfXcpX2zZS4U6YecQLlI63B+GNntwHwZ54adij559eGIzE0vxOVJJg
d56SGuJRNbG8dZ9HeVlj8bGsYBCTrIa3z+wL3LReBaN+Dt+vm6Z1Yw8DJp2Jf2caxHgwK6kEPlQ3
uTjJzgfOG7KUumlsTqVtvjU0OczAewF8Rqpa/E6VIKTCmHT28MsME9JZ6P8lNhPxWhFsJTVwc3Vf
ZHVb/obK3NqVwlaPgkf2XyZpMCkHmwMKOq0Q+sclsPE0O9ZX+us4N4yY4IY8tx3QCXQj4rP+9tGT
CB5/knwhWbjQ1/7ObjZuL3iUDKs9QU3G2fmdlzn35xDe1A80zFFoBuL8UHtpsKPSQRRPG4sZrV82
77dKfo6yDk6Q/af3qEge+A2YN3XoQ2wMu4if6Q3QpPitiu+LTRdF81QWS9NW6uEZA8PEIJTK5MMR
IWIuYdapVLJN+OiS8ge37xxIcB6BU6NHUI12ufzaJYupLvNiGvQcW0+BiyvSfC6cOJOAg34G2CUO
9RKrN3qkeOgP5KlorzUGYY+l9M2/9Lr/kkajtqfsSaZ5i6NgBid9Ycf1J5HY+T8Qkv+TxM0g93k3
5pLLIYgEHngpd93vLelRuIToteK0IgAFt60ED+9HHrYMAcuptdYoWbUgzvztIMfjAuZvRMCx5pEE
r6LOc5Etm7AhQTffy5vYaatjJzeqkqDiLi33iZfz1DIV+Z/Iv+hbPYfwu6T7nXSqF946laTDT0JC
Q79QnRMpArECzE2uL98m/m90OMOkeWI7zpQ1LQU5YDKRboY6IEyaBw389IwnMX+reNbv6H3/Eb3T
ylUPv0ZtE5rr7rgJlJAmufepTTPHi/UF0MweD5ivZEtL0FnYwbvSxHW3jt+3jd7yMCfJyyNsu/v/
WVGgTrgrMrTYHCWFuVsKaDCSjuu4b+Wpw7+T4fO6HIHlaFeyv8Oq8y/VwKSQdxznaoQQO1D6uNOq
nEZ34HURpxdkqqH1P9RthLy/RflCWyoem9y9R5FW4yFuyTqoyyqLFp9c73EBGneCgILMbeYYVXCB
IE2XqZxw1PtQo86GaY7arpExC99kLf2G/w0l5yMYsfuuFlOQMu0PHIGwfRcazAgKJs5axqC8NyY7
MvCRqFHlznnj4SQhVw0D9GPx5towBx9ivc4ePeloFnqVFxcvphO5fk4kxuVpbuhxoNbp5rc+zTFq
92q/KiVhPgImcagv4/T+DM93JDBUt8wtZ0VyjSuWuCoFYlVdDumIt889KwgTuTOyCsAls3E3LC5H
DL4qqEywaY+mgcewdMe/d097MxVXvIT10qPOyujXYsKNm1Y/OEig8A4CsQ0gKrZ58fmo7C3wG/m4
UlMbnxVbirif2n4m6+PB2xOlg76l3PF99nz0PeYHash1ilmBkhfCMmTbH72MAtjrbTL3B6gi26SU
NuCwr+inM0h73Fo+U3lmbHa1+DV7pZxVOuu/ZJeWm+96S+4a4TIt1K24sl6nX8p1zctqRXA73aJ9
G0gPhTqvR/Y4KgFSX0CifRIgNxSvOlElQ3nD4c+43u4qHgCJTIbCVEinPQFy7mxZUC6791DIceM4
G7Cs6XFgplo7m1hhs+iX4xTjkHC6kwI20DSMPr5gwjGCM3u550tQJa7qpdMuhBy1XRCWposnegrH
Pn/gsTgc6ofOv6hZGqvQ02bqroxtRZ2EstblLUG5+OPqqsPV9QQevL6bPH4/VwqSYqAfSiFQNpzz
1FvyrWsoEJpQ5krxsGU7/qdbC7Av4UIVqPEkEyHeRfMjtCI//nHARarp1DkPcMgR2aWFuQERhFsG
8WwVS8eqehmUTe4+FzaU+RJ8e7P5BFsaK5LJ3NXObFOUbx0L2nFxCMB1qap1WBOU6drgFNKPYUG6
P2KseOVtCqgQU6Ca/G15Ut1IENkkfO5ntC7IlBeJehkKZXeBQ0PHnpjarFiBJoNLmx1/oDGXS5V3
5iAG59+ApR+GqczTJEt/TRx+9SLYrvP05WY9T6ChXpcEzYsYj3mg3w9EFD2pFyoMU+2BrqtzptdL
t3XxKAtVvymVckU0yM2sK+eTf10dAG9oyen5IhStrxcrS4D824kKI7yPl56oXrNR3nAPBu+QcgTE
dp1TW0S84T0Q493gt+m+W/8DkNHCbEPBmQH3p8BQ9Fiz0aZ37ct2P4lyo3vIXnmLFRkLjBY1mVAD
g0GGGEpd55AGUpY5uyq/wtPTUzgfKn0defgBvC3lFxjjQgpMRnCkz6IEfu3sYrAZm+zP1FpJ29uK
6nuq9UGe1J8DtnKGcJapCpwapoQW/LfLrtDo0YGOqXezlkk8CSbbB9/blw8hWrVW6qVhJCRf4+H6
/mpHJdbYYbGPH0b812cWAsg0R1kctwq229zgOkpDA6eahgX15p2F8cFgpYQ9aukdFiUelKhaBoF0
0lP9PtbMYo3bQ1+e0RK5VZ5bNlTs9pMSvR+K1QE4aJXqOnROnPGUrprYcFWEXgl6L0RRzOVrjW8d
NtohEjIILNCGEITHPLoVqxWLqUIaY3wghD7Hn9jUTensaYv4DLHtdSZWguB2eIUcdaelg1JPYHPc
3YZJM7ob3tzWYoNa4v/6Tm2OwtYkM0duM5LEnwe5PA1gvIA/E1TfvJ+P+kfXqjhBEKwjfUAP5U35
WT5xdh68ViVvFsxSesgORTI/uT5XHM8zc95+ysVvbQQAGlnSQxF0DX6HC7uj7JypgJELXvMDVH4b
gbQoYazIZlSeduzZrixjR0Lmm9Etvv7DgWNZ7bxHrEPr/heITlSnxlmbDHQCYWGcxR+7WeH27r6m
5kYPfmFLYo56OmESNzvppTmhiKzW7Q6pC7XH9Xr7K2MZeAJL9J/H2aTQFhmjwZKVCGsQeVltTT9c
5HaMq0V0Bf8UFshey2IQx0Qn+KE93dRDGZRcybNAdwu7lcyTaYZ0tQCg/1AGwuyNSY96cf5NTHoV
v8rlcx9ZEwFr7JIVKAezeOWSGJjkmrIytlnwhzQ2rJdL0w/fDvVsZjBE6iLCjSE+02OoJ24aXi6C
bVi0zrXl7wiPOXrW4uf81W6C8CZW7sGvgPOYVWL1rGb9Jfa8cxGrDBwPL8HZl/6PiO9QV43XPf8f
JA7BqeJh1ddONVQWvp34/2vKWsTXPdCWRyWscgggibo6f1Np4JCacU68HPSrvNo7MR7L8SUjzUJU
kxCduyVYylLUhr84rG/+TCvBGN5bPfRLMDOR6BuvMbotfFa1M0/n20JhEKI8Rek6T1aBvcwp+biu
77dBmpjO5WlRfhVhCQVoawdVfT1X1Yl0l5XfBgsfTKCDp41ndAhcHdAnl3vt1miU4V22+dZ8+vg7
FX6Su+osmYWyAR8hiYsGeN4E1m0R6q0UyKgrjN+bALUlAnIRO26eoNIKNQ26+/VYuDkjqNRlf62r
eHI6WugldK20q3f3M693CpMjZljUcBSuNtHvychIg6WWfgeZdyjBJ7tKvfX0+U067Fsslhv7KeSb
PkG6nlVGptj/XZEfNvVSJ3rmvovE+mXjrmShQ0XFOPZPRR08HTl/pN4iV0Xw28JjkeS5V6dw56yA
LPWG3y3UeNurKz/lzkXE82tgho/KN7E02wM0+3GTwp97YgArPHEr53xUwpIcUkxePvYeUzSMZDrX
lWh68kj9xvGdLLcjZ/A0TzkgCG7vPS0IQ1kncy6+s5Zricwdg2KRdl9QdWtetH9H3kxweHw1upUr
AhCFEMt5YQlJZs1/B79J66XQhw+9STAuvA3c5P5oJthfCvzVuDEO1Z0zr7RvaK8B+zeVybwfx8B+
e8UIIWGAeb/YyxNWq5XixN7SYwwbaxXU2HNWQVSzRsRV5vJyYm5Ra8VOGVTneJzpr0KKRwQAQ+CJ
c0qeOxoTlgKpGqSehATVnZUm36cS0XdxqVQIolmvjy/0f+WCoMMd3by9diQ5OWwsIu6NrfpGLa0i
khga9RIGPw16WjwOXZadZzU1H7YF6ot3KWsLO5oh4OYm5EhIex/m+SDU9JPZlKIVTCoQYDtRTxqm
6se1Hp9z4+LOCMknWZSVnOmiAQAIqhq0fhVgnY8Z6xRe2xcHnZfR150vL3pbSh4W4R6mVLDbiF1V
qFs9us7u12CHuL/gH3g6H6l1nm0HuItSWlux0hveW9fERjmDKvUUFbBjwnpl6CE5qQwg9pRWatEu
tA5ynp+acAyMpB4XPfftoh761aYeakdWvWkMkFbQJ0ZV7KvrBDkGtN7/8J5L8Bi25Rm/KKnyqEIn
EKjnTDQv8nxNJuhgFzNDT6vGb+8aoIDjktUqo3mS145z59ng03bOU2/STV7G8rbnq/zr6c6cw10J
U2TvDxU3apgV9wtS/magCxzidK6EsBUChseb3Pf4fenMIy8IrdHeXkP3TkHtf4jhZl+8hoikum2y
PHVlK0n9PC5FG3J/XT8mzc+ZSXTlYUjM3/GZJ22Bs2KkWp7UIhufs0jLYSVaSxcxhqRgwJr8AuXN
YoFN2e16X/fbH4uromthiNMGs7XtVHk8N7Pkq1KsRX97z670/yQqkPAoMMsr9cXejKYf7fyqsQIA
hSaqDP9y6wbDTKm0d+u/4zhqrWfYCrMA4NmM3yRouunigE+aye0kA6054BX/xX1uystDsUgcv0ke
G6E2WV6hFWlSKF0JkUtb7LBKDEz4UBF6nxx7Q96UoebSSh2t5USYPZtRijmIN5KFNirjjrnLJ2zv
dk39TOlyCv77gTcIIgS/b8fETaWS1RyhhY5JnxAgI7EWVOVJWemrT424/3rapfnnkv4wK07LWTdh
QbPa5FijCwdm8VLa5VtnFBp17AJOC9lQoK6/P2CJfD8gPwFF2p+kqRMfBZ1hH+nTWWrYOYtofJQ2
4V6HcmL5N1Mo3pKTJwCBgPbBWGLFfrNF7XfjCSgYDtkCBQxiaNwuDEili8tyBYY3WjYgXGavzSUZ
bV+sjPW6LdBCbQXT9i4zztersag90wercVDgiNjdTNQKrYSBPqgI+zteNqUmhWjUcqrTi7OZkkha
Fl33rICmNwsxTOhek+kGyA9U08HducRd2xVSxkWCh2cPlozld42yZX4DL9NU58EZskXYR3S+1hLW
1VE+wZuML1gCT6Der0N7xipfdv4Gpso8BDkSof0lZ2KZOkNB1HB+XwCsgQXzMdGNh8dhJpIHiwqk
nSTTj3OfRLLacVKqpCDC2UeDnHujJKzaTLbiMOibbqsw8ZSE9El/YuqbWxQX8KKeOEfgx5XEOvSX
+pLK2PmkMeZc06pNF5dTk9Mdxuq+u/JHfiT0CL8oNDZe/8G/+fBbUT68CbkGTnH+63KyREIu1qOB
rse4eSNlNYyX2p25W9aFJsDGSUa56I1e+TA/MGYFMlN2zRcNUlhI7mYZ76lRqgvbOc6lJ7mKUaVf
yeUUtltswvdwLT9SrQg1PoKWs588moinhRYAGZJxMstMKiHdEIqMgpzb9lenEvxh/iPu40v5OQrT
tWE+k3TJ9FB1ljwdYiilVTd9M/5pRG/bqRiImMgDAN5kOPgsQjdv+tWfeLyDitRFSX9XfCL5MXQp
59Hm+DabIal7Ay9yYI0Na+BHPe81PzzVmZG+jBcV3Xla4TNc7y0THX6r1FUWVyjDnPj3V4U1WWx8
aCzzF81o42PJVjrqCia7TUB9j35ygWpZNw+DJNgkdT8iZbP2o5jrCUuY14NpOTY+Hmmf8TUhJXOj
gFWsVvf+7hDob+iO3Pbp8twUDBDvag9vd58wS5kmCKlzbnVofEHZz3IXRInJf93U0IxdZrRakF4Y
92pc9UyE34wZ3hEzDptilhCUgCvdHKPtj/Uti9x89/EQOCtnAzsP9eZqodeEn0N+Pdg5CrYQX6M1
Yp6x1GiHiI25ZlRwFDdGUYXbn8HtThxt96H+pQ/pAPv8QZdKtOEhjOv0rpbjIzPyIeSj5UN489nf
AqmhSBhE7+Dvua5BQZCJsNe1zzjuH9TqfQSsHZzZ3f3ngL1k+7Rk3lPamARarL6TSVcFScl1C/Oq
garFqZjGmNeTjp7yZmrY4dCtdPREHNVF2PloDFsiZRmdJ/+EdpIqvIMpeK5BVD1XuEHt0X/EE1OB
r60YSqbPm2vgYUqL2qtzQZz6DdA/4T1b/IQluplt50+3pBWICkDAHyMU6fcrc8nnfbAh0m0Yzcui
WPWCqJZYGACr65he1uqMOnLSivUR1T5A0iIwHBrtLHcL+okP2cO0zKhId78smfUMt5r0jjf3PP68
I/UdAX2PBD+7KVELdxle94rEzi0nyu21JWxdki39KqHgSAQQjRn5XSN0Hgcf/Uz7IcdNCzJH0O78
F3uSE49/jy5sG2yi0fHmT+dWzbzXAVFvGzM97BRaKp0X8b8MUtDhh0Wyi2ud5XYwjeD96QGABXGC
w5mIwqk+5qIIuJbfVyAKi2/RLdLbVB/mdgb4ZvcmpkTCMbc0etgI67AsunLnRfclVmJjZM82A6w8
1OSTihkUMILADvxh626eGiyvpf5lKzGqj3Ne4j3W4O+ocnzOfqZgLHqMG3vGKKpEp5Pm/vXmuKh7
FDSFAwQ0rqvxOUqPwnau8m7TcsU5B8hVadPM3F6KqObeiuUJjDu877CXvmjrd18fvnnrdVd66WIc
ITOeAFOBq8+Gu0jB9kLPvEms2XY8X5QR8AtrPIKSxroQHDHTDZ1J1rhapzX1+BwGODMWHs7Igjwj
60NJzv+/hVkSbLngjPXX6KQDkmjiCR91e10Q0zvH1foD5wp+iHceEX7Vr55tN74jb9v9urH6A7xd
Xxy1GOohxpJMbkERDDDxHjp7jLDqUQelJeZZk2usXYsynYlm/kJyTC5XssEBuJ/7RAv28IBUttcr
IFeqSDXMZ68NbnKF8xkOJ4jDXE0/7HU6LGo46+KdJC7SytPlxb803vJ5M0SnNxUSJ0IngplzYFI4
rQVyhR5kXSAWnRkVaN6yL5yfIxi/Qe5fFOjCx7+Rh3TnLucWEvzwGg3Wtwuy5gmbreLtb1lqThbd
KFSGWKT2lYbDply8kwAb2GCwrNEvkP1DKm9Tw3swpfeHFTwu8jGKJwxF+d7CBllA5luZP1KvuIrI
6AHestHJM7IgaSuCmnz2RdpRNOPbsFUNpghCuPx/rOSFOMP///lT9myYWojvSyPjL4iXXFcUKRrE
iXmJ7+UGaW5BrP5ACx0w4wwOQZUtaBkyV3mmA4RsYdFXpp1bk0rN5djXenhnL2Tk6d1xncz6WIxd
Jjc9GhtaUJ4Gkb4TX7vJNGUYOi2nB+C1zBE9M3NS/Y4lGZ/UA29ZUqJVWHLhZxVqpinOX3DPq+Zo
WwvCyNyUoa5Lbe4yZM25wLG6IuNIttE3OtHuhaC4X/nbohFEv5jHP1C+Bg1E9yxjk/pri6UH9lRF
uaGaNLn8aXk+F/F7nsFwTqCyn93l7ctM5TYkfD1dBk5yKAu2gL5+n4np9hbBd+1aSs3cM13sSfcm
Q2vwWDJZymE1wBFKQbJ9OZLDPdrAgz7BoelwA48yJFFaEnIAv9p7kWK25aSdHFhahFnu8t8buZ5e
z+zWu+rDUTBQFrk/u1ndv5FoTfWOyhnrlTevM64UBuF+ppYuKgV/g7hMiRu4DNPyivJPU0oKF4io
v6OaAbLzmdQbOwLJbsXBD47QDBrbRNAfmFTP0zHrAY5LFCCJMNP0MprpUW+EgwQP7Yk7vv/gwCbz
gPl16YXrUWa6P3hJRe0v0LyIgU0hygA3JAVgfke/bJ3XQ7dICbOXFsgQVd+JKWC6F8czb+GA1ZCv
+DJoiOqctICgqpKF9jrOka0O8YxNjoMQCQx8NhtKm/ZYFkPC9hP/yfckO/xqHyXZWXziOa1QazRb
XCEfAj2Fc4Ipf8L/+YBK+caUI96yMFEHIG/r9Ew/1zfgnqGiOa41NGaZjIZUk3Dfisa65Lm9585I
eUlRkv0IGOdvPGC2BxNDE44IGxFqHGZgLbakyxk4ArL46beoDucAiDgkyArmJfII0IDefARLy9cc
H/Ms8i2SthscCFX8rh0Nu3LwUot6Py8kJkMpubLtHW9cwbP4WG7TSY7d7Gh+CYt4tas8Hqd+Q4pR
jrt0mjIduRDYsQZ+bXdFYbFz9BBQZk2SbVCdCH4GGDianKqbPU+K2+MC5yrST+qf5OGycml5ysZk
3ryzas1/EiauuqTFNOhVfbMnzvqlAzVAuow4kPO6R2v6Auc+OeUKOpxtDOa+YsyrAvKbJIobAdzn
zXXXmTIWHOZAhASdA55uyMVZEQsMsUcROAkTD9bCux/gHMfoNxwg6SInTLFIsW2P/OYVu+LjtyY3
AhY37VW+KTD8f3M+CNtxmq0ZNkPLvDhxI1THEf2Re35JsG/mhHn2KmYwTQXrBYlLHMOypQK8l1kK
5aYcGeBpxYWd5hedsPWqHp85HET1r3A0k5O8yMW+Sm/2FfeQGzsRQd1LeVv/veWfVlJLgoO62Rpr
kHCjkmaUnjez8UvxyY0hkLhGoAnzYfwWxtaNai/fpnCvR9YvAwQXch7MFtEN4RKiAqeorZlj7Lhd
vMj5MLTKoa5ksgTeTAwFP2CVXPrOujRl7QjTlUhreOhI6Ou7G6+qR5X/7d7HBgNeosgz0o0Jl/7p
hH25T8fsBsnHp0NRw7za5lpAxcJn4xFfMMCFMtCok2k4mPMJTnmZ6Q69FZ7OLavJIRD/lK3qAXKX
8zbv4W4Ca8X7EVQWHfXBWYjSXVJ718gNqw/lk0QjlXsQRsaDAUZqtFPfUkZ8tW9f+WzeSfaka2br
/rasYG6Zt/neXcd7YrteqLxZeBB5CPUE/TJnPsLw8WKCP5nBuPuHzYB/3xBkbPg4TrWzXKl+HKFr
eJMVbAv58BMz73MOiY3C4/SZfML4AmCujAtVGFwndCi+o3g/RPUv2yrHQ41reZlySwNvONbgbs+m
Ic8Foagr/UzKM38agaSaM73u1Osd/qVf8AQ8XkuLCSXzSIZya6glu8YlxtAzGHPLU8OmGUzIhLWi
EYdT00mGjpME7xvsXChdYKO2Mejgs0yjMAlpfAolgL3RkBg5fhikYeU8M32AFwhcDu7jplYUjzMr
Ni+ia7QPRLuJC173dwMfv8jSeLPhO/013ZQJcxkbzhCypW7ElSA4jWdZOgfFRZircrlAJRScGsEz
TDnKQiH9ukIvj4r5QKrmyyA6bKqrMSre3FqcUOPjKoVC99zvphC2Uluh4HjktyQGjhXqRtbhoO9f
bw3XUdMDSIEBtpZcT6Xx8RFeUNuJK1T2/G5X+k82pguYCZLLkHzaMPMUJ9ug847ifio9SAIe52c6
XjmyFSA+iOdtIApHLN4b8+3frVrVzzZrh6FuuZsz3v9KWZdjJA3hEZUwazO8mSzFfwrmL0LtxVAn
hjt7HO39iD6i+D+E/HtV4CGCW6T4XpMJkEt4YMWuv7a6hSUGhYw4m1QK4/0FhS60s+hC35VUfA7p
mVwf+uhHI/nFMht3howRf1AkVOse63l/l1fhGWNClHqb+Ls/wtdz814Dh/yjkVKU1MBdnX+nBbm+
XQ8gXlhjDVR50AazEqOANWRcvHA0oy+0Bium4CYmRc3mJmcZzb86O0YZqOJyFweagb+ZQ41YmuCB
1KWqbfQi6Vp4eXQiytV2a08oOuoRKHNqjVu2Dd/Gb89MQcLWMyJBjrtfDYg0SeADWvCekCQjN6Ex
TTiXmnrHQfG/7xHrFa0nYHooOdB4BUfHDYiPOBTvqaBFOEFg4idlvkqVe5/1Nved6yxefOFsLlOg
gQDN93FBsEQFiw+vwIoyKauVKDkOk15H9uKSCwMPs0hvs7jeCt9w2Kzt0bLgKzSlFRZeSltVr6yD
G+1sRY5oPh1CpX41ENqLMACRpY3NdgWMr6Jrp8RiRTcH8+/h4fb8fSBvvjDzUbxbl2Rp5V3hI8rI
CR0PmmTYDb0EaYifgWxI4qGfwPvvVbGdLgrE9fzMadhFNJ4C3EWjlxD9irz+EzP9yNoSfSMvBJw/
pb/NbBDwQTwEHwiuBM+Ag9vHM9Au3Bm3nlpVraXrTEFh8qD4KVjOmmV7+G6vXgm9viPIISlOGThG
INEuVVTBiKeVPiRHDsAC8lNphUkebxpoeykYPL3ixSb6sUOXllOfHBsReVQ/xfDw4qmL9y2iB8Bi
dYswkMF0HRKHlmc3WKj+Dkw3cq8rFgl1+7L9Y0Hnxom6Gkrjmw0G0Lztx+qqaGzZ0HW57anOXt5f
zmurLsxbrUYrjfkVnHryM6/5e1Pu7A/EIV3KwP5nYnSFRmdbSzm+EfPkrB+mpEtr6g+2/Ip/Algh
b2J+ry2dt1ixJ/OZnJfNt+yT9m9Eb+Rk+y7i6KKfRJiTaHkNvJA8Fk1snrU5capd4CJlPg3vcsOr
EPs3J9PjE47oYkvPvw4KyWFv5SsvvqeljJ90HY4FV+FI5lKNZ2iq+SbGR/r7fEapL/8GwfOLiA3I
KQtkonNMvMf5mxQFV3//5AXD1UZgApSglyk89R23d3JfMsnqKYKQ9y2hZYjcSxRuN+KSoQHX2zay
VFaRA/vdHGFO9YYH4NujfJGFHLBzjReLnM2Kc08G7UR9n/xg7+vy+DHWiXVW0JhGkUouj9rzjPd2
g9S/CNjYUmriur65iZzvWjxRCepu9C1Ba7vChfStnCTAIt1q0ZOPQKOuPy73keqAaboV9K2BtWTj
DOES3USy1l7NsVec4rZWHOMN/p9LMbSerte12icRqVc9nP+TiCHck7IQYzLKU3yOaIn7ZZZayvAs
zCaqCuz0y+zDyFdXLB4Fk03wQSK6In75fgxD5qZdMB6CBtNBVz3fizN6lPIsel3Ix15H99M4mRSk
59H5Vkp+ypjZMdy7Aolxzpel5CA8+h+FrqwypmPpDcs0v2i+UZ2rBDdUL4XOHju/lo3UMf81XcJK
TVaXYqoQRJnl2BCVFfzVGvfs2mTc8TAM/29IqB6478tCQKXTvTKukVMmCo4Q/CKFNuI+9sxMrOuO
a9qmOP+x7JcN6xRaHC/lgI1gAHc8AI24mPvlattrBZswAlYDRhGt1e5yZhMwhrRvL9ixvHy5TJyd
dCFHaQyrohYwP3vRR9DhFNddAAwrDemK39HaPpaunBSs+X6W08Fvg3yB/AkqN+mZQorb+A1UjdkY
QmpaaHziPd+sjKW74oAWb7V7vzPlkqeKQE/wFlYdbHh9uAA68IBR93Ve1HFN/BLQMlJkD2fiKIEI
+xnza3Tur0ozOC/qOOzSfxGC9OThOkcxAo+XcFNJMSq/3GJDNM670QvsmtdwZfK2gPCw5K9JnZvf
ny5CHfdR/VHAk6GbeQkk815fOISWVD62WKVhKUwTt5n4ooW0dJfZo0edRB8GFlSmpnCEFsGohXwi
PKCC+CzKM13uFtswB5pqj38bowR47HqCi5x7u/ya3uTyaw0IlsqDM3piTJLqCfwwhtHPY0t/J4PJ
aspDVkr5WXCRxHb5SFu39MqTORt4y3W/9AUETgoCbxkb7FPBd7QYt8myHYLcGc2xUzMJwdqPbh2d
BluO8TapnCMWotEdGJmIml28/f5hM0W3oNPs/qSSYlvW7b1QZuDjV/Ley+wH6I7vm8U2Pnmyembq
SzeuwdrwMAkqhD8pSnQXaXqaAqkqeAYgFR6E7c9jOwlY5MtLgKpGkU0WUgqbnWnSx0K+thaGbuQM
v93UrrYuoPRFe3MmSBReMZRP5NWpH4r0QO4eDKrZhlj1IMt9EIgjdtC9AbDtHV2jFJcjx/I8OYuG
fZ+RVXTk9iqZTGIo+OZ5Kr8jKHow+IkPHkCFAwU4l8k0x+dq1evmjvOBb+0JtsI4exOcua3+m6aK
PztVfGNheO9gLv+WzPqKdgIA/q1IwNBB50+FBsAijPZWufQzcNB214Ra2MAq0LYUxTxck4LWVgwV
+z8g52qg9SK+FOexW2SQ8mRO9L7LSr9kkFdod8tTyTH5X+nfOWnfHdrUMECeuWzryc7O3o1c7IYZ
Hn9TKLKfTxgDhWQXVUk68J3qAsx+27lKkx3S67VgLBW/GMBrq5zEsNYcNiFkoObIU8iJSMVOrZCT
zEDUTcp8jtu0EDqd2AP2cRIUkCzK/AaKdEN8FB5CKHNO/QPe7sUozANVbQ9cl/4rJbb/tH6tyEFm
xq8I/4pOv6/FJyo4aNqXaMzm/CCyAB/3/7N+D/RN0bi3LfsfQKoE0/+gLusz9d/BgjgVN5ON+p8y
A/hbbJ6vwnCqWvFqK2B6iXi4p0rDrnarTPMkAB8xKVydLMhZXDDCOAsbZ0SJULXSSW9gvBaNPnZk
JHRf9TaqBJ4KQ+JPmRVLgvA2z3QFeqHeMvev6Zm5GKjBnSshY7hfdRNvm43MtS+ZBb6fXI4/733a
isH7/S7wXjB1mM6J5Hn6Wr2rAfPrzJAQNNjSZYT2N+ToPgvEJ7+BtoTpA+1aAOIcvgfLN2Ahwh3s
Kt61cIELGPOF4jVHQSEr7lIkol6N+iwU0UFZoJmQrkTaRdS7C+Qw0fwUW/I+o/jpK5DbNkXS3BkS
yIs+E0mDsrpnNWN9dNeRrvBRE3jYJQTVd8P8+5nKUQnzgq+4uXeoBE9L95EFcwRiL5ir/EnVXGkD
KLGiTSzUofKL1tB9x15xgHrTC+MMHwzxXE5PN6DxeTXiKwOoawpDjq3N8d6Td43wHU/irsjbYm+s
8cNUP1G0L7rF6rBAlpHacbVJqQUsE2Y4ODZwoEWxhg8uaR8EcmEQK5VjY7vMbKgaJ5wfjE6fm1Ho
8lUfEJhmKo3GWPCVf3p+rFSOWBGGs89acPgPkcajYQAWFtA7s00gFSMEJNpaMND4441GA8Vb3jZi
qLI0DKXVCw56KcsC/+qN/xBNvqdjEPn5Cue97y9ZxpQ73fMA2HYfwvZ0csUcV887vGtshyeKlF7h
f8BBY+XPNlWRuy9kzgN/sxv29H/4PigVy3eUY7rjWrlxepwYaNj1rKuYG9JmurKROyvOm/xEiKD9
k8YXX2AyBUEOrd6Plke9Lij171f59LyrtmuX77bECkYv23BcZJ+Dw4xtpDHAmPWPNwq59ej/3fi8
Hw0JuievTpBvhbJIHH+lGSrD8SH8rEAJJw/9EbqDKAXJHRW6kVjfcLPcGo0XCsL3aBOfk9Zd43IN
FQ5p+z4XTqfycuvMmmyyNb6CsbHSoPo3vXCGSUx/wvLQpOshQKPAPdubbTKYUJ5aqRv3QTWGsfPv
sunvZfRuNFwCN6WxBjSaLOwDZFX03lv9rA7ulQYDdfc/r4eOnsfw5etxlo9pNyVkTkXStKCwNmMg
W5zM+L1sHCSxbWZeI26TnjrqDK7D7ls+0xu8xIhZAl9jGm0QkuzFVTbKfJSRxGTeJOcHWQy7Awl5
kHgqJH4cRZ1ioB5syWd7MRSFwcqYBrnGV+HvAdXJL4CwX76+Np9dZx4cQ9lJ58swtrrllhf6CAdx
45HRkCwKvvfn5CLX9awWsuyBOZ8mx7mnSO9UytcAUfqNu9cs/L8qvbjkuMVlLKV0KTTOrdRI1Hdw
NQBp10z9LfPNE1/eVESr01tkgAc4ZX2KcpD8kdL/1but5LUXxHd8Rd4psO7PZAXYcUYaggPp8au/
d7bmS4GOXt25c5KPgHy1dBsptKZmbGXUNPfVmbArR9JgxkS8G0M7JjMg34jnh2/L5oaj0oJOzoAT
MjNI6Lu02c9g9+if/YelVxmEfz+Jh7eSIvc5UFS7KS7v+ilAeDNmDjTuaGo6uQ/1QBXLFVtWhiKL
QNpvOrk1I25JDNjxa+1OKuO//V1PBzBD/pAh2hJY/E1yNPgMGU9UgjIJ3lzwJagu6NkYF3bHDYnP
TKBlu7pFkbZbaTtTCrrY05k6/Awa3G+hC69wLu+UNxuXwPdvZQgbOQiBjeqROt3wWjRjePk0JLlZ
I9WtZWgLsfv4VbAXWs7pDAE22zv80inrudTIM+I12bf6JHj4MGY6jvY/Y6mtx+X2v3IDj0ZIbvJl
oShOwtUAWMavd6mB+SKTghpm5FZzgl9zWCofmOhAWLy6PhwEP18H0kgC3xLwEiPrYzYyl1YCzkf7
G6u9qYSIr+w4Gf8kZnVL1EjZfgJHhu3JHAkd5RC/KHnonWRHFVzAXGvI0gjf4uxAAVvmW4vpD+6H
I36857SEiTzkZke8yQkANMGnt8/8YhIjrgDfeGgO8BnLCDT+Gbp++78u+C7p61Y515feRCoOX3ql
/MXX2lE2i7ik4w+Pxlkb0Oq76tQWQvig42mQVeWNrtGLVMR5LK28HCXwR8OsfKcTC3RUZdHsza7f
zx3wyUcPIu/HeDeXm/AG0SkamK2ryPpZ0vfaV92uIkE73EjX6N0RfgO1DBhx6kEBECImCQp605UL
b2pWJdi3L94M7u44bLLD03i0C71PfBbePIQP1G9tGo0RoSlg/fUtchWW9DtmpWqAcp36lSRdQPyn
+4cCCl/5KbmajwHv3+j+PCnqZSNOQAy5M26Z+aqEt+Vi9SW7ngfx0KdaZY1/FZQzF0DydYhcIfNO
8xwBHTkD2FpDT4LGqt+JbeElNG0ZziHSvgbXcKfqhuYCcam/+1Pl2bPixx+nRVdyCb+3VocxkoM6
6Pmv5Xi3bb4h7jsP+LOobrp1+ZR20r4BK8O3gQBkrR+0qfHsYTJWq969p8Kq2x4JtVwy8zP/gHrk
7BS41Mh8V7s2M4sKSizr+nJGct2dRQwRTpDGdYh75yfVjtTi0Rh4EB8QiNJ8YH4rMRex4dJZ9Pp/
7PmES7GIe//Yv33Gv7HmhBU+C+LoGDIQh30R3J0K4aJwP04gT9B5zBnoLzGoXmSPHZlTu1txTkq2
bnL+ssrW3/fj9men5+PTwlJA59FYux0nptxSHvA5p/+SEa3shK+h1A3nvjAaZMoaZ31l5NTma8dd
7XsFHi0+7ovuwS8VMFpD1F/pQpl8AWXyNW9OnuQb1gP+2bgzPlHSOUV8Qqne2fIlS8wxOrI5OdlJ
uPgin36XgaludWSzhw1XkfhpaDDv9nAlOdW9VIkkzuf62b4Vz2gzcSe6Qi5jsslt6q7EfCippli9
mChlYvZt781HyCGc6WiELBqCdUxCgG5XCvP9WYv5Xgj9Q6igruzyIdEwVBOPSJWHHEnihnDkv03+
S9e7wXk1JKgnhLF3hsUFbCnlzm3trW9Rz7ZcsSyT7Imv8nXCxrvu331DXneK/Mr+60XjbcLNR5jS
RST5xzFmD3w0qd3bAtvt+z0OxmAvyR3LlTb8gE4gNg+dWYukdaHnjZ/OOeqAd70S2MhEfSn/g5w6
A0f5/pkGtL1eLLRuWtidPWTV1w5CkcELL1WpDDd0MNLjG4ln+IGFfDz2460ZyWPLZiytdercYxKk
OcrtNqf1ySMGN98rRZHojfY1A8gFjbGpJNoaf/13Rgmcp9zDZ7mF3GY6j9AWVKaPL8LIV6Yz1S1A
pJ8QMwbAILbh0ZnjPYjs4PRLmWCKHHUDStdR2gJv190yehUDi/ZxPRS1nJCJiWwnsKloNZyH57Cp
q3xkQDAAmlgbYKVToJH1Dc5QWeCUubJYD6CSI8ei22luLZZV/T7XKKaR9UcMHDbmYgJ9frnKrG6S
KqIW+9zW2jCPQy/Pe+kBYXjbAG2KPYT1GztR8wKC3syhMF/DqmwTj+RdsdLGYa8S3QFQ5g1rLDvp
2V+Jr78aVTZY1EZ9lUCNAH7XVarpPCL2kZ8hThUGp9B0PWUM/JZQS1VYJCr4ML7PW4BcmB5limD4
zKZrQKJ3/rV3JzRWX5NLpPAKNEGwKe3SsKoJDrA+zE7HtzmXVMz/Lz0rR6P+48aWWP8FUpUX5LPE
EurnNvEK/5L099WEM2DMkZdIpFexjgkto/DJKVrXYmwXEY4kmT5z6rslEMgXZVgfzy40sX9y3h1V
Up6VBnPedTyxM0XAUm5VqdCCmjmGtUTlkzlPTg+p7UBQqBFEhu5SzHOFPYc04gD48sS5bu2w89ZK
cLpW7mUnJ5DZbFCWbSrF86LcRpd/Ui8cltG4LelGHBzF5oVlASPbFlmaRvv60Bkz87iGO58GPWOd
/FPV7FxHC8svJ2spK9TuDMs+foiQRS5sdX9ezdYZj6OBWUOowM6XfAZ+q9yO0BWa+rUHbPz4ToDR
ioCVSqHdGxI3c1OJYQ5OCB2JHqrl52BVo0AcOyN5fh+ToIxeahN4ryw3I11GBXcYX9WxyOINLU7w
Yh7aloF3AcNtkCX1WGHxuBTeoRY/j9BTueh7VJu2vTQOU38Zj7pMy7kXP/ftk9TygimIfNEZJ8kD
5uPAU06pzM52Sd/rAOssidB5SlMOJrsB1kDrrOzZepcuZ/OUDfPrK9GVHidE4qKJFX+B0LM6idMc
vsbFcuaYT1YT/XIhsEWa9KXI/0tCZAoCKA1KaaH8LNJTkyIDTmdTXKiyvBdLEF6Qwqin6LAXeIhN
LYxTeHB6FJU3NPnQY2kN9P8UxtszmJ5sk+/iww7qiaDBK/XEnQ1nlfZ8oGPimEC8vyzb6ueNIvi/
LqYvgvoU/qtQzR7kv8USZVGgN5Cf6TM+1nn+9NkNTLRBPUv3vUD0UAo/3t4sdFsfM21lK5dFZ8uy
TyNLSS18X1hZydA3pToKL2qTKwz8QK8TPIC5N0I1Txv5TUHgt5GwHJ5m6zZCvTMd6HgZjONov1wF
SFBqiKiISVW4W+jyXQZ8UVooq9KUyXK6F46EzSIPFTR207avBdHrbccc2dz5MEQkrbQrt5XpgZ1x
uViMuxxdlvr+kR5ln+1IDjMDi7eV9QXk/sWNHQ+Gbua29mYP+ghY/m/c1EfANP5tfxrU4vO+xIOa
U3QdcE9ZPuDVTa1LD3oZkdOfe2jezzhxr+IfeuwFkXIVsJJT4b8neUWosQH4KX2q2u/WUDzbeam3
A+PAK0yWqi71AfiSGQ7b4FWR6X7q+oQYtyOtT1AX6aG+sVqxsZVeZE/VluuZyOjalUnJkXGeOBRa
5jUi96g9w2MBEPltrteAvVP10m9M6Gl8oblixvhc6U0Aw4kIfeSpZ4xglPvDpv2NjlAbiiemDSg4
2oAVqt/jO1sZsiSw5ea80wVzIWMmAQplZuGhyM8WgKKnmUTLsQ+R2LnNFk7jticvs+En3Q+DmXNQ
Cfb47xpxxp81hr2fFj6NvdKFLBq5GTK8ddgy5+P3YvgdxK5sffkKVGKoOEc+xW5MTe1j3XrLziJj
J+9SXkWMcsEwniYHHuv3pJ2mmzosP5cW5psgrgOZS+aQrz3vJjRjTkN6enZZHsQnUkFYudXR5fKj
f/MjxczOQzdGS8JNVFuN7LJCp0Imobpvrz9MwCUdDVDriLsHOyHMhP0Y99ykpq89+uxklCZ67154
xbZf90DM3bZ2Bufr5OAJ1cL5SsgLyMmgS3UM9M4nosgQ+AKlpdfTifh7KySTERL3tGBCTzxMG+IN
pOvu/ATH7EWpsVqxLgcDORPknPEZJ/A2ORgg4ia6xZaATx7U6S2TxYK3zoq1K/5fGrVeQFHy7AZe
pwrHfrBkXeTK0PTHOv6tI/NXY7a8gbpNwHhkPm6mLo/28vQSkDz5rYTxPVoGHHblo558G+a9R1RD
+sksQl+FWUlA+vIrmmyiZH2KZEBMM8hOiWxU+2vm5mILlWjmuRY+d6WCsHayr8RHxYwF3Kz0bpMt
tT+5JpbYTfzQ132XoWU947w6yQKiVhbFEUM23J0uXJLrXSRM2/7b1ULl1oUDlblH1ueSiDjl33PX
E6NPzkF//Zc5I6im+hr8GEPMnQv4uJGe8MfMN1hYZHyeIGN41Hb6ZCz1J/vYLmXfGKwzrFlCDRIm
sbiTKYnFHQo7Xh51A4GHa0kVgFme1e7TNRDWi+iDsfNBFUtfh9ZjTG7rWOeib8ByC1iqsTkcWPTD
MwqTgiK1Wnpo58eAqwIc+7DgbvnVrHrWXCvzRM4Inj1dv0BZ6+sAku/VHblP2+Kosz9hltsBgok2
8wlrC46VnmRK9/11PqZUnRhQbc8SiWThPKUalZTnYxD/loBwii3YKWjcAVZSq6Aj8iR7SZLNzAJn
i3T3F7jRxqAiqpZn5BFzS5Uu1dEEH6nXLbXAi4eWCBKHkUo7ag0RR+V0akzd9jK4l6Sp1MZmUqhU
hRfcjWYb+ntLSnBscLP6cRu0jUwTylK8DT57S91RoQA1iX4U+ES/2yPDXK+5YwreyJDo9wTbmBQQ
QgHxPfcKgr+FTtaqGwxfGq4TRg2hPE8jgH+aTAt0wPa1xVcvaTZijVjQWNgMca7A6OI6fg2UsKS/
ghBYyicBsfF5zDakFzziOw/qnYARLHef8V9LRnq4FkbFVxpkVRaYqHcbkrJuqRsFB1mpLvTUZPzh
7ENe56AhShmi5/HJzuT7MrrweauHZQUXq7h1jMYd513Jv3QZ92vlwDMGLaOSk16BeRAG/dUCVCxG
CBzMAkwEqlYAfFB2x/kHVMSs8goDzVo2PL40w5bWq8+nTILQ5YQoJktRKPoib5fQXnck8Dllk5hb
k2NHOrHSciWvvuqMPF+3Zy9B+SiNWGGCO60vADa9uL6EUF1VGtDyFYti9rq3ZpIOzj7+e16Wrjg7
TIfQPVKm+ZdY6af/hphazeeIEXxrXElrNhuyR0uKrb93u077r0ioIz5iWOn/7AguYWaF9C9dsx8C
9EKsYjXTV8Wi1xh6m/lN4FOiSMyJHakZSFmdcfyhK6Vhu1t/2m7c6XHTNlZom6xvDr26mJX2uDOA
9fNwlWydBzqyYxV/9z0foHeiKAMDi4cBJgucs+hL8C9ImYs9mAPQx4CClX8fjVJ+KGNU/1MWBslh
sCkEReYs4xf8EcbyrYnAIm+r2zQ3QzBfnnuyfmRqUk0nFW4H1rsp7xMt/Tbe/WR/Lt9o9yA+Tvwi
Ths4VbGwWsV1YICSw1Gck8doXX1riK9uf/3NRvPfodjSFhxDuJQtKO3aV3W2aeOmwoyvUDtGseHx
eOggnBKD1uTBK75GTT0nU3F/e4H0Pf0hNreGRAtxn8D+ubn4a4aH0ApEc0S2SlhKx8EWrdcGrTTf
4crvCpO9x7qG6cjAM8AEomKafz37Hn8aCCSDT6FLoqw/Q/emJhKaoYszCJN95K+cS6olIWil5e3k
huMcpEwR7IBcc0YfpIFhZdrf+shyXGsKK8Hj3cTBlKqJOa30dsMD0Ppp/s7arkiDPel54Ai5OcVN
z8OW7jey+yMsIYwq0QBDJ3eAHaDOeRAZ+QBtZbzyaBGK3c1Wr6eXcU909N4BqvzesyUAlvkAyi25
0NJE37kkfDWgEuy36XKVivwn9GBRPqd8NcVqtbv3cYey5Zxl8Uq7d+SuTWaGje+mkKLUXuRhB0fu
DvEMnZT/AtdcG4gSktfGDYKy91iDUBSfI1JMYgc9QJpgz4BJ9akJpUrxG2HldQlIQSelo1BvQjLf
3rKRtf6W8SHgDj3GpEGcg9DQti4WWekQkHHIyM079mjhjNvUBom6vfuLH5qiCSGwNMCKEZn8hQ6R
Red7fwisUvNbByM706SHlaQbdz2ZgleEa+stEox40BR25/GEzB5lCFIGfJwkUOcr8jknjS1NvYtn
n4CE357lPCI+QRhsa+fx5B4ghQuDpkEVKp4/4iST93mzjEXcuerRTAR8Al4mYbhZCddjP6NVRhHz
ERoWh5p+yL8DSGc4KlmF04n88/hCZF5FKSg6QBOToDZ1LYOy7pkRMovF39DqRpIs2F2EBTJ1V5CQ
SNy6dYbS2D/tZKMc5NohK1IGJoRGLamPmPAAqAJo6/+17O1/EV5K2v5fQqS4uR1atGYTC9MxZc/R
Eq+5GnsEYG+FWYPtsJvSjZDOP3Hb16Z0ZygWiqJ5UyiNE+1MMfl18BiUAhpb2ikkku3igQ+QBBIx
0Ac1IBMxFsV1XrSZjOLFTXMGStIiiSu1/hVznxvsxQgt6AWPtEZltaO7mVcqD1GVj2IpUBYJopTF
AbqXBOFg3uDiUR1jrzGVHOlbSdDwRPA0jbjq7CWmwO1Ovc02XBJ+hwm1SOZGVmJvN/AgPeK3JAL2
gVUbnYNzBF5+ZBPSk1u2i3MdsY7z6ZgaCYDhS+HBtO/M0xkWVS+DBtZAvljGBVNlDizz6mPC+bwL
X7F9hfgSFEWqDGwxyJ0vdF+IaGimzIl0f3dvs8c5JTz6lmhjhi/CDkAYb4kSi4vwkJXpprXDSV/U
apM/5UedKxhnflqib/2BXhP+sifekT34Nxj+EGBsw7kTSsARb4WqWYxPYM3t635NTPNLca92Lhta
yJO7BJETVWonXFpwFuEvwxIpG+m1p9+VglxxRWj4iYqaIamrVRIeOdDDpN6NUjJoE9R5ivKPYjoJ
7iBbmaKGLYzSBxk9tKDLCZswznyud3PyC9Dw2kE2Nt/GGRuZt8FhL5I1ZoQ72xwrcQUK3jgGCkIw
eiHwgjAKVfzL+lMRCoQJ46M8JbOKBeVErg9jKBCdh87LAE+IaPBVJNuoC2dWUjjvnsBSyUL/aAiO
OOKyBWoYlGHTCchBpvDJy+SjOn2iC6UjC9oUvJGxsgnRFvzxnUUpUbUo9saiBqSQ30EJXKNEbEVW
E8p1PcIFzniVm2ueJl3ght671eRLMJqiNdaLUg5Jefpn5hhca5Mr4zLXOMJF1PBTvzW+jtwB2m4A
X8/oqFzJTf9LcrlBjLYAbF2tO7Sf7HiCakJFcLRzwSUHtlLbOudSKYzQjAFyTVncPf16L4L8y68Q
kZM511RY8LDVOdfwsEirdqbXMzRz7T4AJF1Tkd5rcKXE2KjJzt9+FRypIp1K95A0JYx9UiRg4kF9
nfRimHIt4oV4S2yOpK6ZfBaT3O611AZfEhdfjgvl/1ClqcU1jyMlRMgw7Q5r8oVyCoLXpKJ+xtrv
cHStDurdx6hLGopI5sWrY9fW4rQfbNWl0jforPrFqRMKRYBQ8za5urGU6x74ueAXWWkONCRrfYXj
HG8NKzDJsfr0JKcvf8kihTJt88sZIh16uArxcVAVrxAThSWq8369jzIHyXHDzke62uFt7kZY/EY3
qA/ySIQo+6a4KJSDe0gwI3wrCW7E/R7m7RqaVtQWMm2gOBorWlzoa8UhRTpyW5gTckJtDql9LVIM
UBUZVbmzF/2k84jrJcLDepEfajYsFzMKzRMx3T9PKtTHJlGFDn7IDK7T2D/oxfFy5ryGGmVe3Fev
Lo+wDXoNGcD8LnIKmn2o9qyDFGMBxHWvhKK+4gDi2P9I96ZO9CRrXqqTjsJzuc5YGiL/PmF/3hGX
qRn2QnX4eCNO35PdKKxfat3odO9Tqml18ZwGlSuH1PpWYstE0ID2BsNqRRer5EqwfRpN5BdmeGOf
Ztux5w4pE0jlKlBn7QLRNouNuBxMaZN/Cjbp96plsCsNG7cVLbRjgAOLPjaBKutag/HwB/x0Rn46
ORKCxW+HuAeGS7LqVOBhId6ddaFZuczUgUUvP0PdusMmAcwPAMADO7hloqX9+jrBhktttJaSF//E
5PuxrdluwT2pmWYNRiHwpvsS3HfxurYZpMfJIkC91pRa48x1Q8/6dj4vglMg6KP9PjT9yTlg7ZSC
gMV45wSIlozIOzk6cEGHFdSDJstkjuv+WijwKaqEl/dlj3AHX7Tm8dyAnvP03OQg8Jz4EIOyha7z
FdxJoxMGHh9Q4+Ol/5HNwFArzI4+joN4SYCbC8z6+yarZHRdwCJlw/S2Y6z3T6URkGt3Xy/0W6Eo
fssuq2VEdg4uISCRmWWgekrPoba0eDlOSVpz6dhGKXqLVjDaDVPVffGx7j3/8gHT314QnM810ijT
F+qjykaypswjNNmtBM1A9Y26A6c0lID6no9YKH2l+eXKkmB81RaK0/pG0Om3VPck5/aDXJos+yF+
wCyEvMl/Nx4WO5S/2fuezwe0lOfVZZPwV5WEtMz5WHTUoW0jB2BJgRdOBCbaq/dQjApB9K9weDlM
m/8Bu5UEFQ1B7qhrDPqrSy9V4gC+E1eq2kq1cGJMBy3O2cFu5Zogym1lDhxdVf6Px9/NWMpEDYV5
Nsm3bER4g/eHoQHXfS7aWth5Qiwsh1rz8O5tAvRLdYu8ySXEXiIZrtSGrQ83LM/OynlSAMYTzRsD
60lbGJMkjyf2SalFwQTRI7DzC30qBfdbvBmlURm60SgcfoVaq97mGlYsnpIGj67zPZH5nNJc08P5
KCBBthGCTS405JZFHc0mk+84MjzT5eULOGf4BGFYr3aQHEirak99/Uc3A/kM5zV22UXQMiu66QNm
hc9RkpMlMAzEWFIHpaSUTG/skaetZGcG8fMLuXnzgZluxN6AGEw6W2Hmd9s/LSWh+uk5HC4vJZ46
lqspmu7N2j8Dov7MLNq+3sosEJBd62zMuZXWCfptLOKbnAqW2KJqjeFmhQwl2hqcyT2yyASDJeLF
/moMndGhmEKaF1D8K6+XNAergh3ZMg1tfSHmbXuBG5C0gxfYl48BobKQX8dAmg8fZ60lYsTohFRC
Mpb8dDQ6/URWfnLmcpRQSiv5KJjqT9mc8tm/Z9aJdRXaopElKYlqu2uqoRFaQ5dqKkYAtJ8jGDWT
3ra6vtDL0MioEktrY0L9pVsl71drLSqNv7MaLHsGrhyHe7L92T4hqqjFKP1TgM6DX+J0E6o+hkUX
VXEwP/xSwh6wV/fEWQjQAE+brcWidDgtiUqaxs8ZOtDyRK/FPgzAUej4UlxYrq2rkb2H0WdC9pvW
T9J/5Y9x+z9ZnJa1Pp87oCWJkUiH3V3MbxMboQ9IXu1r1uBRPZz42bUzMlfpOeQ4oNyOMbIZruhi
QkAlsRzYGHDx0125YmfGK8nmm5vkqsp1S5jrl19ng37wgQgY0VqBq4lbP+vl/5TXoe4U9bxhJ6HA
sOUU1ML0FN2q/bpUMUSPrY1CYpUu4FeyHqGqdIstiBNGyN7L9LIY9W6G66oDd4EgqjNLCG4hO/fk
0gIZucBmy/DRUHEWG2DVeCiYYaBj6pkWYjWoovZur1wywCG4nmMqv18ETkZVPs6tlIOEFiU1ui7T
/deiLI2DXCHiAGJdJqMMvpdRZjSwXiOeYbrRIsBs0QQ6Ha+M9f/QsItwGjaERXSxatMIsF1uQOye
Q6U3T4AHzpbrO2xYYGr2twLFIpcybPpWXYD4y7I0On3zsYjIQ3Gk7e1bZYWWnHmlHyXZbSV4CFVM
PVbFaWPd//vaRgRua/Hd0/daJWKosTDwJ2Kpyk/vdmKYF0Lgu5+x4DIfW622xsqW03pfPQWTC6jc
TCy95j6dcXguAQPtvCxyUDL6wFQXs3kDJRIccc9Q3057eYitHBWgw0avb9yz7Sbz6ck+NvgC3mJd
vKT3WhbgQZ+0Z89JrVVdy4SJKwZhHzfKvQI426J1AxsdyNs0rC78kk31ZVsZ4oMtAqK+3KP4gfyJ
MJbAXpxg8eMrDrFWEeznFCo+n6rn/bl9LwRNOye8+gWXwDlGXkwW+rgE8h++SwFrMMNeb21adv4b
UYrwlOxkEV593VLwFqUNQu6xf/K08Kp5HhxgeMi9gA+TWKyqnu5DWq9IgiS7Pkfn7pl10qPNL/Qp
ZQ0wz529yfS1hDcXXo69leNSCZJcavLW1EZVtPOAdbp4zrOjSUMs1u+8H4sksJJTV5k5egpVOPcX
AbQfG9Sz4jDnOiVHQszyxMiytQjDMEBfTLHfTe2oORTw2j3v56wXz8yQuqa8lE16L63binTEwmhQ
7rOYIOpo3tpGX791czg6hgsgkZs57GcjRxTv5dQact6xtol8jFdQowicA6yKbIzvBn1u7i+IKDkN
eI/SL0awnQtAuAR8d1KAM2vlrbzm4VdRwj+BaJLskJphIVjNF3CtcAAItR7T5YtRkG9l24jbCSq6
SoJQzYMTHWUPzVPyfsFXp1lFu81+Ut1e1lJKqfJ5GS6tt8634FzinljZViNTMpnkfalEPRqH7dnD
ek9tWMcpTfQO+zHuG73Koopf6hQL02z57wX90mqNPs7PyONZAz9PsWcwXym6n9bpvmKoGk7BCw33
ryCNbiHqQc1dKy4o5eO7R59Omn7Apo7F7An2ODtH5JSVEBObzBaYolHjaSVdjF4AD+lnwTVzQ/ll
6WSR3IGPEHOJgYkuQCKWfsqpihmH3IYqZCEB1iOAYR2FDythiU/5zoStOnrs73BMWXsOzP0HqzoF
x3HThWXpt6ECBP0BcsAqFc8u73cG/CyM8bZIl1IgmCb6rDI68WpJpMunwwa3Ng3abWc0jhJ4H91M
5wDeTBAnGfEbUN7nI63DD3ImKXGsNptrloQ/Gge9s0WQJGmzcbWAkY2AcOWkAp1VQ+S0SnvuenUI
+FwxgHNZwj5s7jcX4ia5M1xfvCMlSP1VppCM4OrypE2H5VJa8TAbqpepWC0tWqtoV5DvvMTMW1fp
DqDA7rWmXQrRUHZnwEZ8poTMafsap40gwSvs+5X628fpl2YCSih6y4urP4baQy78zVyM32bKeOYO
3nWRowg8oGLjrYgmlrz/gYTzAWZhWwAL6VIFj9eW5JGovvRRGgqax5ZUy2bxec8Ip88ufoWeA2CJ
XXtWrIi40bGnsBSIP6zFVYUl/Ut5+8w1OY9aTegShz8RCbLAAYF3ZRpqJ/7r2Nd1+cPMRBiFW5Fc
kRGMA6ST9W90dYWjvOF/sOk9ZvBT5xR7rFF7021wm0V1fauRoXnYxe0IhJGMzDxvO6Kvd5DLJZFi
o17Rh3APSUIkLdPhSxyGoNmsMy3UWr7UhoiVnhS7wA/0jpKkfzyq1GjQ7IQt9ftsGU2iqc1GA2ui
wYolBsgUiAUjQoOwzEwmQkT8yts5DNTmRor5VqGFBjvsIlHkOr3r0gE7l4hOx3YEnpzUq5to6lJW
4lC6WjFIDWdLYoozJ4OYGeu6YLYTebSA7SQ1oU7A1HWRfYwEPWTLVg3AwH5WiN1XJ09DJMGxn6sm
wXcLX8zAT2Swf5s5ioJATlKdAfiNwKNvVBz4vSg09mjEqZ4XrYkk7fjA3Lqdx+t/hcLLVyZsyzlN
dPwDY8LWqfVPokvvxSBy7NkcE4dZzbt5YsEsjq2GGYE4XubU773AvBb85S7jdhaPNGqCaIrtCqoe
YWEmt0/Vry/suH4O30bY5la/49IWLwbPl/iSdpCz27ohmx3hVcoWqEcyxivZgIkbagj2DAWHXp0y
e5pMidQwXJ+Mq9n/HXXWrMJdy1ybZSTG4ffNo7BaZ8n0sg+/pWAwz1+TzRGJKhHHmTHSATiK1MGW
icsv8WZRMEtHWRkJR1NDXEVgIq0owRdrlqLL2u+SfDvACJTnqmXsNkm143KnVMe4wwnGUnH0FEMQ
54gYUhQ5tJy4NQ4mhsfouve+gAZTiqn7KXccdwHOeCyY7uOunRjmmKaxoHHf81bLuNydnN93t2Pb
398HfkUECag6IhFbOcuuCihESOecQu+zaaZ2ILZZQ3ujnmnE5Kddec6XQFjPX9TsRcdjLHN6KsNq
wQh6mdPgsPJ/0rT9PqntZGeSoBmUGrzkyf5pk+Vg2/CaEQFdMkv49LdZvUBQy7KJr2RIJTk7Wn94
SvFTss79MAPLDC5WLqvpFbfZph3xbSnNgLmBJe5dW3CL32YqJ4CdziRi1uBLNB5r0/dY/IlBIcEj
qjLrSKWGgT5y8PHfPVCPyw9ffc8UHCClreJ2nD4lnRQliy+W/4n+FWJs/CrIgoEub7JvnjHjaRxj
tVZLF9S0hdWxkouoncsAsilZFmhwj6si9Oh0B1L0vJwq4aPjUdcQ3Y2V8Zng+yRVWUeaBcKxfxf5
WdBqxGFwypFC1o8HaiwvzabIIQbd3muiel46qldIZG+nxShnG7bSt1MBEwNf6ZbiCtRDr4JpXjkU
DPUMg/9fxeYrwZhA67jNuC54wC2WS1zJFbOwDpml2dC8B9KG0YLn6z6JudNEiPVfVWIVw5dIyA5x
xWgjEPi69sxg59k72RTB2h6NbWRjmIVrzGvbKpn1MSvDef9ps7Lpr6moMSvdox02ZgwUNu9drh4L
V0rAWtuKjeTT3aUS/3hPvPMdTH+NGoTieJfvcz+hFPogT7VKfSZfi3k0m9CnbWNkId3sCU6uS8k5
QJHV0tOQr5vs35kHqgBuRW2NfHdGZobi9iRbwWlDf1B2EurNZnD9rpVsb+Tw6MrJBYWPvns3p+Qg
roiw4lHCph+dvJZM5p2AcMh1tQdn7O2PwflFPLJkldxsnJJak7+SJVxqKIIt6eJ6OwVuzp0ZEN6J
6FJqns1Lu6W7h1IsLhsPPM1Qio1MWgN1GGMcXuhVQ/RKSHY1B9JE1eyRgmlQo01F3RNOsogpwh3U
CwgfWenqcSpTTbEx0ZVnzCCxW7MAU1AHATKPGyIXWx4hfSR2LKf/tT+weCoofJLHViaV38kwb9Uh
imonoXw+jAX32VpVGjXE0HI3dGO73zzal2/F2D1Q9Rp3xI/2s4MnfYe+tW1uiR+rdax5R6e/tx7q
cD5G4gjyfk32UfknebFRaXVzXDGA6aNyioXqzgJj9HPgGTm/qTJNU/oasxUYG7g2kTgGEL3Qx8Ty
YRPw1fcyattZFau/bf3YbIMjIsSOs7pjSybyYwjwcqooNtmZmYS0cW+CtSojJw61suSKBcVb3O3T
Aal7ldL5jHdO6EhGptc7Fb4V8HcAG2c/ah1C8nY3xsqeC5hNCg2srktKEo51qNr3gBumuPAn+hl3
jh04Zb9uyfeGOJ+oOPobrvJ+t6HilsO4SoRwlXIiZFTeyyOPhV/XFEidPw2pI0UwBVoShJLAuq/X
yDZOmQZnrY2MqJ/mGrDqJiI2U8HMdTjzIbF7hJkVOQrP+KgkeF1K8csiqza5CKGjfetdhjG5YEwg
cajoNrA86DgBZNf6mxsopZ5A7qTB8gaajBOQe3SmvkPHbHmd6bp6Nkdh/bsdrXsfiQGAKx7mHSMw
i+RRa/YFH/YXwpSKtwxsRJdx/MZfhqCNBw3RLb43lLmb9eQD5fybCB5bzfDKojb371oW0c3gAVIZ
tnQ1EbdJizeXxMGetcXovScTU8jeCwYtTpDXd0kgopDqdvJxkMGXGfoWzl41PgLqzXMVd8xOnyR4
vP7vR6mWG0UsAtV9RtYgS7HTSVYDyC+DVMlhjn8m+2rdRGt+qvLxUcEcY9v6MDvLV1jisGSLtxld
w1U/JaQMGiMUYzUZE+QDUfnhv838x4u5AfO1mS5EXK3LpB+WhqFyTyuZExk0GJ5w6vC+T8Uxrzpa
Fqa9jwdEu8xCM1csSaxddsRORfgQCHtwr8vRal5ZR/ZhwuQ4UQLVCBM4QDXIaa2M5bUAJsLaDnEq
mrxQVyiXzc+zM7e4/hT5/ZKzEPevI4CXj4q5FdAkVeoGYatJDtxU1PKdg+j8EAgFBh6JrRon1wr8
9wuouTYN1MFed6L7fKP03zMHl/T4kyR40BTeoTWhgfukvio5pVL6uD/JcndN9ndxkRPPcwfnWwKn
LxjiIvOy8AUweaGmebhUs0/OhVHg1jY4CCzXyf/NQaX0lk/DcrLxwt3WrEDClX5zziz659QngkjO
TDtcIaoomp/OGNERP2I4VfRZfPywgF+6zgDcwZGoFuGDj3y6Ga9rf4V7zQPiO6AepTeyc79wimSb
J3lNK6Bwz8RCitOmuBIeINDEPxEVmhoYwzqH5LedScbj8HGzs8HU6izJdYZrDqSSzoY0O3SnTUEm
l9aX5S0YUWezWOWKoxRBFqZk2coJIELbYLSADiFUb82HVeWyC71DWd1kyHjaBnpNC70ftro7+TGF
IrDSnOmfFNgdNn6+DyyQi5ShYwujXlOy0olZBkhxX5NdwrOJPzJ0Sr0SHqdcU+XMv2zXLcxM+roo
dwLOK1kyv9UX8MdAjK0gIvrX+L4qnrbDi4Y7XfmkzfT2ihVYSnHEymIZpU8eXfypOuMooV8YweP3
BNbgDUFkkhBXtiTzfQxIF698YXVcupQ3jOjgqIVs4M+1kwmbExrlEPlv3N4OJgxl2sGYEiPK5s6p
GsNMucDoTeaH7pT5r7Pkvkp/e+RvNV1x0bBhxHzEoXyEjU+uJlml1+dsDX8DVxtfBgGL9VgkaFsS
ElB/YZt4S5ZMr/XW2DTdPMbYj60jrOsao0BtGGE7hPmqFJTmiyBmbObR2lRwFcE0k+wRgyJAMNRi
WVbivQ2msf2vEPQ+rayfTxrLJTf27id6cNSqTQNze+a6/XcRjgJp6KBdL/ijGZxVPXsoXDMGDiQJ
thlpVG4U5GQ9pdGzJFJ0iy0ApoAl72+K+y7CDn0+NyV17D9n32dais5s4ORTECcSxassMV1k7OgZ
P6K49k4X1zQwWiYfSlrVaMn3nZbdHolE1GAHMrKdcp8oXqfhDUdXR06Q6Us9ik3i3oyxAVmSlqCw
gR+mJ3zfjYgUmHOQcP4V6Zjpt7hCm335Q59Als1ggG6EOP04eub92KcEq3rkNW1W2MEihqI2QqLG
gZJvAEjAcrbfa8vsNXZRZyC7l418uQH2X+wWEb/l60ydnFeMKfjEFBdhS9LAsyt6SJd4nmJKNRSW
tboufRBfulZ3lob7Rl3bP0tu1Jf080MySbxsqNcZHzR//iIrbXhchACya1fX8TYLFOUqdUOQyL9v
m5cX7OLtLE6gtCqJZkHdb1r2SHmOwuXhPg8k0aSNcWxDQDgJDm9ZNJXhrbNM2Ni7wy1lrWrWQ/KF
Ny00fhDDUFhtnilZIb6KaeZvn8R3S/xsfZ2HQQLkDQjo0QHMUc1xxnxsDDsrtZxIBeZh76MM2DYc
+kJSrVzOf+WwnUr9m8Rn8yo/EkI3tc8NaVSrvboa3A/eH1cwr73SVM8mUjo2Ns2G0Jp89pxNzTda
Kf1tJ0/l2GuPSNDNCYqzJNB9NpqCLpxdWpILIRN1zrt4SizgzHycXT6VgAx4XePnSjDVRv7omqkM
+vw9N2Nc58WdMUFawaAe0VK5Vsg0vKS/3plsVdgJSIdc9F+uhXLLv9fmJHMs7zD1gY2gKc7FsySx
mlmjI4JjkZF1mm3yy8zMjS/2+CQ5vGKmTbVfoPMiEwdjm7/UbY2iJ1AKXnVwa3BSo1bgjCAzgxE6
31YfdfSNovYqnm9Qd7uJUSyLNf+AHGQpscIubySZEdBWp/RrLKqRUXWP32mq5YdWiYCCVjZoJYVb
55Z8DhaJBug487q7eQqn3ROTzlc/0OxabEWvKhrAC6oiiksDMhk/3zr5AAfcSRCc0buq5mL32Jko
fOEzNaFp3dtfvonygXRHqQr0tDOi+BgtAEXICaXVDR131+4KRjI+eDoiUA+XvjSsVbpX9TPdGOub
EnauEe4f7e9ae4hVNzah7F8M2K48oUTzzzPk5Mmtqh6WKnlpvhNS1NQAEGRlQ/bmvwQvGkNgorEo
jg4qIPC9lR1SGROd3MXiU5ZrIOos8QjydZuAKy0gPqe9yjLL1/ogWpTp5AEMDxVMNzwHKPA7xaPi
GyLJJp1fClueV6BtDL9QnCSO6l1J4aiCzOf08P8SK3IQccxW9fx10FXKG/rE4zErWFg+iotywkFZ
d+4HhUOXh4Id51ZiWp+0fsuKwxcJswb+6jGW44qFN9xB/Okdc1kyL148qzKxbKgT2J3hPDQt+N/e
fVSbNyHjJ0JsfiDWxA2wcStlEYsmh12Z942gbkWoIAWzqXR+n281JTYuDasphAsEC2gcpbpDYRC8
yAUWoZfr9s9HEx4EyLTVzkSRanGTWpbEmig+p5V+03KEsQafBfm4qjEnDYMshaiTDQD+FXWloXtC
IrLrBfv5AL3/h7GNTFAWsk6yI6dsgC4tnnKnyTGVcBHan2Vd/y2XETmjC3kPlQZ4/qm9QttX6VJV
m7XXVqGYBAxoqiRR+DaUt8p91xWr4q8hHpBu004w4hhcf0NpM/+UbalcV6OZY2H1qgeCnG/3Ms2V
3ltzzJuyb9HBozVjmqHap5BIWJ3K09wxueaYKLbLcIigb6oF8NMaMyzH/8hphf4hLEdv641EmR0M
LpCkpB7pXKsm5f0yM06CFCBVxkrEezngsPsaXbyzGQqZFRZKfE5Xy49yXG1pDP0ytG61Ik8YQe3U
JJPyRYXTbxFZurxOgdQWB8uCzhpYJEEPnpA4KMsOcfM6PcSIbKvzXIGdirOxCWmKia+18uAqqJ+2
Rh2T8OrQTIfhH7SZZcreQJtVHm1iPsyGPgSdqCjX4lMNwILOXDFdlQLCSKJBInivmN4eLFzNhSHx
QcsryIFPezZqya+kAZsv/DUetJsMpQq9SZknNYsgPd8NffAMK8Z52JGkAAM3z+cgIRzH44sA7RVP
Fuz/PRPp8f637rGu7CnhykxfGwRVIYQ7iZ1bZbTDJXTA1pivdYsWFbnHGtOcGrB7TsHcyk/P2z27
SXfh78vYT+/D6Xl9/JjSoFOXs7rFMRz+dHMM7TrkUrecdvO1VVOBa603FEjH7OZN6V1dOcE6IFca
SMbRtymAA5ebrBRuexQiomEWRjGLMU9A2Y51Adlx6rQnGpgVqtRqKTCM0h4CR0dvVj9dDnCy4OkA
gQeFIvBplDcWPX/GEcZmPnyg+R+pSWhNgo1wX6gx0KsysqEp1ZfbiB28PsVVAnoCFs7kOviSa3ot
CtKyzKnDFyXAZfQ2a8uPgLt3fsDbpA3bZI98EfwU8xDQDkbCzwelQfDoQJaivpN9ZV7YHEiSU6my
KRWQZmORdvmuGX+5WAwYi83Eea5YgcSWxtTkWjOPj9Z5k6EWUE4JrGIpBjnGS59bz6yYTMtISUKY
jweIo9gW64P+Hl4o+iXFukUPD9xf526Aoy60c5tgP62b/nmswJLhYckLJSu6Bf13E6xs4u6h/MO/
VTIktlRJPng/pQW7Gb/cYTI6MnKRyUI3Yt4d4123QHIxH1XgPALIjpPwRraALg2kfy5MYBAzJkmR
VBj5Eu1tWBW96Smr+PG365x8m+Hdw1oHeupP26lqaevVn/MyoM70yi1Xj2WxCQJf+JlsAGRdjs5r
ZfKtDyRQ8iQe21JmdO8Rm+OpFm58wtfq4BAhMc5jEl6CzDnPQT+qXBFHyMx2w+YYl4TtyEOjKkZ8
584v2ottN3h1pz6baFwH7L3WtmspRwkZXiyZwl0+MluOIOhFbCjEDvSwOaWiPT0+L59iQI/1HgzX
rv8koqN/m2l4i7zYISNDyTOTZSMSm7AcMan/Ol7zSN8RkG993ZSf/f5d/iC6xVZHIHPTuqCCLJWR
jxabh+Lj1iv3s8GaGPPFk/WNjwxdkcHfaMgn72fpKoKMVxGJmhoTMIl6JZ5G8PzyBeyzwKS1vnzS
UdqeQKEhYQ2JkGxVUUbRyplTWXTeQl7OXJJzuG36hI9Yfa9q7Waa49hzuhnbzbAedA2f8HARdzHP
CwIk8ECcL7XUyHXOv/5LESzbN4gjXbmf36aeDa4BkJIjGv3pw0OL8XgTlzZzHpJRZsxJx6DNSoVu
MVm28KvqI4Axhyv9GxVC6cRu3aN5lRRcfOhNHXtN/rxPvCGEJGn1jHCHE/w6ddnf+TEXtJCBQwnE
jPCDAw8Kqt86VP94GJ/9PdvZXGA6vQZDyLo6eoTepTkkYs0tyXCQwibSc5uFICxK1T2pkGqth5a2
N60jCHgCbsULAMw6OXqFBwbzN+0G8gRv7g0C9ISsJrv9zVMYVf5gEohtHCoIC0o/MpzfQGdBtIms
cHdmYEMwijtx2Or2oB15YPoHjnUqoqU84N/cTdGyUDlfib35XaAx/ZvEOY9wC0pklcrEoB4o5FST
MNPIf06+NfZoM4CtawQ1WNZhXQ5hSoObrcJOalbRTXq1bV+yy6a95Xn3zvMrH8Buw1qi+I0ZDL+B
R2lL4UwY32np4Ys+DqgyYdDQU8O7/3fBumhrWh1W4IQdHwluTCuTh6Fi6H+EjSaJNBCpZsCvs0mo
qjUOiJRJ8aRpI1/XngUSWJdYCRwXG6DdJpKh9EHAF2++iwJ+fyIxzchgsxNb6rE1byHV2XRYuGEx
2l32TsNitmg+oQlGTdNO73Y5Vo3PXTUC0pWwofFsVuZgZzIRimbjV8rcYli8jQinuIgNdwRGlYYX
MJqZaIhfeRH7pVeuzJYc1QEPrBxF2bzWeqmdo7TLITzttnSq2QvfrE2hmwFOmytMaVtp3s4UvbOg
XE077EMfKjG64dWBxhE/yjWCvoaPTqHQnj5F0HFqzBxuNqxuMggjiMa2ZdIisJVNsxV4Op0K4bxY
0oBJvu+CLa0zLPXXyCNnRyvf6TAbU/dhHUjIxlgmZbVswZ6HWhdCb6spyCMjFfYYFDEXtQyPmqqW
3zJSQkV4TOg+rPOOAkpYV8nD5zDQzeHvHe4AAxRRkVO+uBRVU0Znzhdxwgc28sWCjWxIlBPFziG6
HP9mAI1gr669Se5/G3jfPNCI5QMuZPnY6nG9Jm2UYaOIJ43Uboz/FzGtmsSuIB8UCUPeW+RQfDOo
KNnFpSZ6ISnINhmGWZ/0QS3LzuiD0iQ6V3IWgIOrNd5J3UmT3tRHA2Ik13yvOLhKEOUMXI4hGJvi
m511YFzXmWA+JpqR0p5kJuTc31j2O51ALDgcCLiinHQpT6Q9KVhZWC0+88evwLdphqYqCjYwnbRa
yeNah++OQEYtGHVfTQ+dSmUsdHGhY3zo5YRJFxkbEJ4Ld/xWFINPFnLIDWBlNCqkBBoZy9oBi+az
HLVf6NoPyrHJu/uYPCZOTUtmK5vPzV9wA2Mlz0/qeSD6oLaDHeUpWvvw0akHBhQL2oJGepthYXAc
nroom7jUq9cRlD/X78ZRiGfxwandYRii05X9u8unqk5n7MyJsm43M2XQGFIm20NKWAO4+22OoJ4E
rpZSdFekSiTmdyS94aSPLOdvClplwT0X375+ZAKoXO8Y2VvA+Vb5o/48TZHE65xUygSNM6tZmcL7
G3zcUYR+KCF1+Gie1ZYIhgj/FMzHSkl9/L1cpELxpFkl9qFhkhvOl/jvjpRo6aWrxZtIhCgIRV42
ZYavIUVbebup+xOr3ctJ3rGygnlMbQJDlrQFJmFDHgDniVg/Xojf/Ug7gFduMa6+jIaNR+sQimrW
98+qRrlxXFSVCJ+9l2tmzaSKEEvdxdL47J5c6ZxIQwBciVucmm+G8hx5PAkfApyhoE4qb1JMAqMT
Sij9QbBh1PFctEu3xLbjPAc+jGB3pDnRNS+LdcekfcNfvNVrtpckqsTn7Jxa+FoaBvYwv0kQmwlQ
hmnoq2L3n+4hUSacHMzxV3RiwE7w0PCwf4xWhktJNjRI/+m59JgS+suTXVB9vGjtCrW1G0FQM+Tj
LyvaNqDKMKT1q94DzEg2OIu+5qKyVMlxjdiT8430OUoZIfrw/4JlIrYB/0G8ynRNuitPoUAAswzN
2XJHAaSX1oCx6WKg3iKsygWtBwqhIZth+Yxbduqv2s7xSUeqF4bpjh2IZjaLYchmraL3W8h2c2k7
7XutpdAhPXpb776QHxcDQMJmjfrRHyDgckYFu7Im32WOPl12arEnP1+deTSAS17ihgU3qt1ire+O
26irC6ZWMsLNC69PBMzK2+wLy/EQ2X9AYTxVUhZPylSHXDokplz9E/c6zfMTbARdrvSJFy8CRpS+
SoqC4x28IDWm0ZtdSkVSIlYMb+JopcLqVO8p/R7EN/LLFAQBkPdX1C3xSuJUTOXhajoy84Ty/gHy
GkPh+jfuwnWZOyi4w6K2lVVQUH7yBtnplvL2z22HUFcLInbDQuMqIzXai2hg0TZnfSpHDkxJSbCP
pQ39s9T1v2TuFYgDL2m459sTBcgkyXCWQqIweFPG0GLlOZSdJXuiq9YtkVJxYyRhgjqtyBQPJV8e
5TChIjbFvGpL8hdfQ9Xfw4tbWTH/8uw7rWiJMI80BUcRew5+VocNQSyCAi5q8B5765f5JVBS4cJ5
E/px89nI4eqTOc/4d7/yldSMlEthEkgS7qwzFR7DFK89JTbFs/Y1R17YN0Ph+f37ZW2QkTefld8S
NzAVM7gYVKcvdRdqaOJbh+7eztmFep8MbH/bZUSjMYclUeAxUkgUEGnjTp1gULLDvVL3nfmR0nPt
FN0dKlOzd3Md8O4cya3nM0OF/cFgz2lBMiJTEinNNLgjGcifcdlrSThsUZ6PHT0btlAXsjraiuXm
BCwdEYpt7UgggYX96nUPe6qw37HRN2Jdodka69dj+v5N2WmT8ECdwqSRi9omjSSX50A/Cyp6qBmD
1IWtGLJad5u6gw7s4H2Et6+vKJKh3+DG5KG/F3i05cSEPuYAlX+0IcL+q1rrlfeokQjYPj6f+qQG
uMw3Gyc3ulr4D9WZ6W1zs3KnZ+CQNdFfGshAdiiVGpdBdDMsHsbJ3IHzpXo+ef78ZB8p0YxOuWGZ
+ou3mWSYyW97ES81A3ZqP5vG71VcsKreYjPFbg7QcOVsmElUUixy986TfQ5mE56aHCcfirpUDVBE
ZIvmKhrFGaI/0yuuBwjVLcSdPij4vzZ49NB20Pir/O7InaS6T/vpBm8WOzdSYczT9aDP5zQ2INGN
A6daK9EVRt89LlO8N6BTXmqab6VyzxWxe0Z4DHYRrE+5OuIT2XZnhvpErWHxKssuGSTHQXvzhJnc
scYkRoXue/1PfYrblS/ndaySyyYTGvx6y0zLbgYVnK/KkY7OD0O6uTSGlFiYgAZewQeySx4zwdoK
5RabfowqIdk+WXe5exp4B9Y+GBMLBWADkjZnq+xla6TLWiufdXsgrsCt2kOYcKyXKo6OoIkQIFIz
0UBSsGNcjLSndN5pyKXZw/bZtpQrO6RW1fDKeB8KY/+JhkJsd89x6YNGcsqeUSGS0+WZ1H2gzTPc
Z9Enrn25Ej3QItJRm52xFuU+AXmwYRV4Cjxe9ww4Jqz8afBtsD2j8r1g55FejBaOpVuNF2LtLbTu
WAh5LugiS4bt3tWPTbNBuKx/M74rtLlT2MfH7xIFHZyYbheWexb96U1vOUfD+mlRVE0MFv5H054r
aRq3r2mVTAclcj+TxV7rXXE8TJQPqxpxq1LU1R3u2Wdc3D/ZjpjuiBXWk1pn/bCsf5EgSuRb5nLT
PT6IAnn7sm0MKC5xvSPk6EwiBgtz+wLSXuASnv8BzomcOJg782PwIzvKYwWYSEpmiPthGFJf4cUS
WqyqLZZT6X1szH+izIveK0py+8bVnqjqvtJ8CCoAAGhnyCKPtWnNCIpD7dnq9OhmtyRDjHMZpQ5k
W7W4VHPzoFJOskuju/ZMDg0Nr5gPH+8StUFbzuQZoWlna0df93UKSHpNJAjFVrREvge7p7HTaNmt
EkYSSgaenADqEnTroKAxr7HLy9xDkBSiUhL60ah1HervAhO0x7mU4Hywu0GQpfRztujXR4gOh/vN
/pZ3aR724h6VUAK879sxH2xtIzgy+fulu0SOqsjlz+I8fYiVcu1blscz0jJ3S3CnzFcgK8y/ybF3
UMcQbEEnjRiMXlv5XZDWjWtTkuRt5AUTJu95sma25/yKVOKyzpyHv1Vb86pvWJhugXjWg9SkOC0u
2YJ3eJOSU53BILEporxuWRep8GrJA0VIauf9mzzPuwS0vPGkk5+6x8QWUFVNU+b+yVzG4dAIxXNh
VbmA/dWVO/9cPoyjwY9WOfCVuGC08Tsd1SPN8mpXpSXs6s4Rwi/euxoK4IgLJeQ0gBrtv9cJcDyd
rsKj9FnJDEditMvskrXWwTHLCZsBUbnnLH9oLhy+tVncTH5qC8Jjagx3+wpXnVjr8gE2tC9dZB6P
Zwi2+Shpd4whUgzMSzpO8cZefdTuXx6Bj0+rCi3oq0KZxsydvEvJmoUupp0ZoDmiW0d5E21Bfkzs
6E8wY751+/rGIRK+pjgx1VtgynYAf1uDSPhR5A0tEjJpsj3y2pHoD7u+nNCY+B0akp4vPlW+fKRK
STe0VVFiU6W6UsLpIFghOHnWOpu9z/h/5pDQ+8PufwdLiIVPrPmJBxLzx0tjiuz6vlzVQNKT7urq
MzdQr2Gv1i8lRK257R8rpG4IQEjbFN/w4vOdl70KZ2SXbOyeA1YnHZ2NuSIssffsr+FH4+W5pC5W
m1V0EbINGCap9Kvuqr7x8S1ptsX0JHmEWOLf4vDaKfSzUM+EApCOdrRbEe0NqrQnZ3TplZ9COKHE
R4b19NxPBHBudvym2m4un1RQgN8qFIyJOAzuqPdI7cNdtD0XdyPB5WATknUm4TXj6jhzv4uAH10Y
s5NXSNJddyUvzPjwNFscLvOk0w6IeqQo/GMExxCPRir4Gc3WViTJgElmSC7uJLMup00hAL7GBe44
SfzshpS/+NxdL6/jNKBs6RXQyzn5KQOucaayshDFksbksQ5ghmrBr0WSsUeCRDnVIfpZ+xUP5n8N
o9J9i23CElVVr+GljOM/0nKYsvskO2hwI2AeKXb42LjhkYGgUAe7y9Jq0kZ6pTYV0eV4LVCSqG2T
xiY1n6FwuSKENq2DjhKW34aPa1kKtylJROZsywwQ1NEf++O6Z03MHUrki6gKPXBF2BND0tVJtoUc
ZM6rsBVB96qIcEN2sO6q7UHl5GSUK9nWMIUAd4aLrdE2L/Q13LEny6Nm+UIA6x+jjftUX/uW173h
Y2bmbnWQiRMI0GEp9SaMC46x5x3N7y+We4ci8+qwrCLC8BCX8knmdOj2Lz4wZQmtr2lstwsSSB+M
JUMB+WBW+LcbgG2uvckCmMs3XwpnGf5A26TNbc56X30BdB7QdmJLRSecexELBY780bb7v4N2Lbwq
SCM4Z53OxYpKGsNlmOBBOjuUbNkzv8I81WamY517TyI2bVWCwJLXMlZS0hJQO5iKYFTIYqKHctT/
AXhxLt8FkM3SThiOIHEPeedwiuAXkOqBR50deiGDgBCe1KA6qx6E4Dqm8pRa+euPKHElPAnukv9C
MatGFgG+0C7LkBZ3xAwwBP9Btz+f7Z7cRQZtipuHkCLGa7nUbjAV+Dfd6T+vjsX/blritgohc2FI
IKLenNBw9cpEuS1R5NfIWzegNpQgBl5UO/LiobTn5qVrT0Tjy1aB+AiJffUDqkJlqNEu64xCJYMl
ayIEgjmx4wkP/XU4wp3N3y8XXsEKYSX4nu8xCtdcmxqb6Kv8tGcP9t0aHwK1r+8UJ2uVVc2roHuZ
KlpXbEb5odFysh4nyjRaYAL3CXG+7Eqlo/wGbcHJI3T5o5bVeMVziEYzxL4CW2gStV1oOkuAHgDn
jacbVm+Ycy+VY1WmktZbj1CmEkrSaRIOH+QwAAb9ZZ4MjJ7HqwhfmC6DX8FnoWmPn6k5HUbR8n6M
BkYW+RXKxsLQqNrY+rCargFDorpQtrDvFoSnEQUJGg2Ts5F0hsn0Q2zl3VQQ2wQ2WO7vsobZM4bD
EMCHBMiwqMG8n59a7pniF0/KNXi+E9URTwlr9XYNVXpRbc85JPt7jP8bxJ+XiazXa+NdYsLctZwV
MXrOeovfNaradN65gp+x2CyjKj9VreKFkmRTlbl6dzcSBRAzZA9XXLo+tjF6Ld2Z1EW6bgpqw363
4dCYnNyUJoTypu9iIzN9uctzIi0Pvbg8EI39dJtP5sABuijtR7VLus16bEmiUvwgcCRKNud3vLFZ
nDUgpFYbzbmuNo2QXiD6kxkhQa6HWB3Xum6IrpkVv/3LLq48gA5rWvEeQ7iKiHFQ8h9yQryVkmzM
x17krdL4r973zyk7rD+6++pnMEX84WZZaWKcLzkNkkOOgOjPgE5E4Bu/fTzaukd8tNjnCtbIhWRX
rw3VysAEJhPO/NI9oVWjkYTrM08PWSOQ+MzvhgV5a9TeMDGnQPhN+6TR+wlyjb3pinpTVx9rsRnn
Xa3R5ieidckBz/4Ig8BmfNwRPjs0WcAXT6e5QGnqBX9QMOVXBsWnjJSj7pG+/WaEJC+hh6VWaMmu
yKYSgEjJYOgvnRWmt3BPFh3I9jrXbR0UVK8y4s+SbuO7xj3TkvfTi8aTzYCwUF1lWbW9pxEfw077
qLYTv6qZ40N47ohswgukqpQqmPq7gQPXfl13wzMZbkjfj6G5HD66nOM6EXetWmiob7McQoZ4KPSc
s59TLZ72+6973kU5zhUmDoctqKpuSwGpp3tB2iWavKs7wy6E1ahIgl4XENgISbAO4aDZQtyHnzZL
5brcKzxjgGYMT/rBoLK4cNdOF5QlPWOncf57a8JMccaGlMBpELw8Fo18XGVGFURoaJVdkCaIa+yc
lU5hOnFWso6DI77yB2JqHGV18604sduareY+z140jXTK84je7Tcam1QrwA/zf1oUPAiL/4YH2/f4
yFNwsm+whMhesTwgyb5iijecp5B0sHcCydoyRna4uyaSUzErqDeHZSwSCb4oZC3bQydXFIMYO1sy
X9LjsVeFE/v4rm6+ir3dwXxLhbaJ6xgjaBk19+t6J+/w67cFLisJPJhw2rjkXOsNwDbb2kZFgnX+
D3H4Q3B5zNKIK6sx/E3+P+W0R0Jv1cphROE+WIxWb34HQBOBOsM/7WHRzSHCN3mlKvZeuxNSLGaV
ZVJKKIED/k2t+RhYjE9Jmcv29x+111ljP2F1mHrhVNH/06eY3NvXYfTFD/AVB3ZgFYZ4fbdsNFLm
SLsDbqMbs6FHr5DCJLcveb+95nIDqwlroU0yHEB/fqIQbAL9csJb2AWzi1lhOCXmF5Mvzy0tGc7A
K6v3j+bUIaT87oE+Lt3hqu0/q6PbkzGrZNKdqHORLYKB8d6u+iE77GPKstPrxeEWoqO+DtjGcwN9
VxWR8O7UWyo4DR0+5k2JQktmc3Y7SqEXdytpHwPc6ntQ9m1k5pf2YoZKad/Thqo8u44WXKKHUBk1
RMnK9E0HDtF7sMBFW/fqXD/ZYepWQvM7Lih95xX/RTK+LYLqxMS4chrYWszZW1Si6R/9ljnxSRSL
oKNuh7gd+TA2TuFiXdJV1U/vjlQqt/ZIfprzMLk2id4l8bdZnBwL62gaVlcci+nyrZxTokYFCBUm
/cfaEXaAP/vS730pykAyptmgZIr7FW/t6vbn8CNLL1cxQ5nMRZvs2XfmR5OpWfmzJG/i++XWLpjH
4bmQPwFaWsCGRzJLIz0cOVqawzbRqMJp1460Wnxkk9j1YFyubam9Vvf9REiMjFlwh+uMaQqfm8CP
HZLOrh7WY+WPkCIlgk9n4VX8hD3y7RhT2mR9X8mnWBUzqESMdQVyk1fz3oS+pJca9TVLQpm6DbcR
htWlOWAfqMbS585jwVtdv+VPQtEqIasWpqUZ9bCzHr7pAzL+UGoxCpS0igpgAeNw2uYXmy6IFo33
/NnCx1a5pfoQbl/agT1nfyQ9W2bKoG11nns7JUOIoD21nVIA+UiM7Tq2fRG1Fw0/MYsbYVproO37
JQRwm/BgxIcvBcBz8yfWf+W1AZX2vgphdvX4sBh9D1xAu6u8SwdZOZrPc//Zp72OC0x6jvQA8CL3
Jk5l2lZdnDkem4pmVfSC+MfNeron4cxVr7rHJbZX43m6PMpEdMtSSVNd4+b4rPWIeRtegna/oBOA
8vJ0caSFmarVA/sk3PYWXFoRNz0WJtmwLa+xRciEBA6bkJI5Gwahu6BH0/x5TgCBzTdmhDcCUqAt
M/SKfCsGWCdOYWL+3ZCRVdFUmfIS+C6evYkVSKi8iJwl4ZjkiX/KRIqzXBzr8/JV6BrvUxfL9IRR
BXz1y1r7bIe3S4SJe3oPbVIVtl8ENWJXVIpKu95sHRiXBwgc5/vElRx7gSlNEL/+L5Q6ZHekWG3X
xXR1iNbt2q4VGvNqt/XBbpsAi8L+n69YjN2Kjxzw4iAfzHQUb31k/AfUa8anRp5TrX5m+3WONoJT
NputDP+zi/NSYJYZ50bJKV/5NS+WoPp/bcvDDDkDK1O9KoN2eNdDVXgGmuEaNi+LDMoKA6Cl+7eZ
Ahfa3nwqPUA9PLtLT0gvUtl9+VUcpQWhGpkHzdymze4IrFfzavKO0eHNA0Vt8Yeu5ke25DBCqAyQ
1y06ptPMK21vAUX4YYNT684bJ5zgqKHW82MO82WLTRKnEAITBPfZPA/huhs5gc8dzqDrWGp76uJY
yD9enudPUX5jzac11gg7qAJTsb+3NvrkDCfSkHvF5h2EGI93pEJntytvHPDi962QODWcpqpuAmrg
ozKCEXdb6zuwK8rANuwkAwNWURiZoiIUM6ZYP9AQq8Ija5n7xxqt6eP3H9Sv2OIMEW2jPhxmKGSX
tVHS+j78WE3NK8A3qnYPiIxbs0FMcxdVcB3kIPdhduxv//shXv/wCXpdm6l6L7PDPTa3gMW7t6/n
TwIgKWu/CM9U+adKSRQGsTrnv5ttmbOfXBvt+H91gbQM9Y/v88+LKASMrxuleG12XNk1mu7/dGm4
hShfcGDSgbu7b66Exf/YRJkqGfLSagtberc/ufM+MP/FanlWVDeDURHBJ6eK2UCauJFqh+oSfKHS
2MzQ/Pur0+YNRycOc4EvA//jI4VkOfM/krQWp+OU5zh9uzZQ8LxYtZmYqlB8jpn2cyl9Yd+w2rGf
nVpds0hnQQRwCbeVcsQt3OjdasXnbnhhbWp7mHpyO2lV93CCdQA3V7lYf0YVq4nnByBMdgVXbW+K
C+fWE1/ONSBKyv9qG7IrWvWdLSuI1puPRHoFsIwi/DhG2gYFwnE3bDv2u2SRS7pllAdATkoFj2rc
mBuN/8C/g1s4GsbST5tRpfrmzX28xwSuadmiMOP99oDoJ09xOfl+LTFMy2iihjbEZ6hnoHV6kQFh
F9YFjlq0wreIMRBLsGEuTH4W2W/WAVM80I6WaT9119dWDcw/f52Y8NrOBBnRAlzi3mR9Cz5lYxBQ
PC4Y60j4ZkHiaE/LM+p4L6GFiy70zZWvPj452TjH//f+mEkcHiXdrhPGHxjmRg7ULUiL5e4n+n+1
SMzkkrlmtr/Y96U8fGAcgESkjAUZXVPz0h77hMrxTevmEDcZwn2zL8LVejliwieO75iVeTVdXPcA
acxCtmtDnVEn5FOphaxBbyrWZLpYMPfkhQptxGxLd5jIrXKbkBCSKBt62kliVihLZICp1a1Q23Dr
xj2w376+KoFsNkg4pOFDTGbrDTWRwcbkqZKCUG/OAKaGiJBADCZTlEJqvamTsdBO4p5oR/u0gEY7
8DMUMkCbmGFZ2JuGkV2hjGiY/kGP2Yc3Wb45RSJok6F1+l4Bpk9fqsmQsdfeFJAjZZyrW0jFwx8d
tcdCUjTXMUuaMcGwd3O6353NuPJqbyCWsSxQuYTAdGMOlbarOy/aLyFtWbaUfq9BoU+XYpOFdq15
A6vVcS4ertV7rL5k8caZnMbVLHlwsREIP1MlyBuNat8Sjqr+HhlCM96Vhr+GyUoCvmO+GtkVVQ5m
jmUkQg4d6rE83Qh6mJG5QQSDtqA2OzPlAYbExWvv2mNiHxa/tNQhxJKObTEHl5M9vVN6ytkLtVQb
9NeRsTwtZR+OlegsjL47F+H9Rfyr5xxMSQcF5qtp9zjMeRPzfQBTEhCZYhpkguaL/kqBjy2Hnnwi
YCeSr0uSszeyzq3zUv+wcj7EuX2B+40PnPPNJVZ8st0iwUPsN0gME2JLaxBirkgK4DoXO0NdiKJf
4piLAQZSIR8ECa4wCAnyiJPsEERbgAVesvhztWbPD5Is7pDxbAeusHm6fnsc6HtoHVNS5B+A6CTl
iCAMd7YwsohvAUgvS96Rddg2gvYkkPIubBA/oNWNn3X/q3HI5A5IGKpPgTH2YwwWQbnV1V+WggCf
bJMA4ngsjuABFtTDGLyoVrCP5e+uVNQCEzGUvLjrwL6xO/Id2eyLRckLHUlefV4dep2UsX9olO9S
j/Ffv4lmmMk8iNo+JNexqY4IxzUFJyGtpe+emmTcgeQ9gdjd1FGVmPULPO2zm7sX9zKyvbzH2i47
euCLl4nQB2cVl/i37gYCyonjbduAWVR4/pQyPteKTT6phuyx1A9UJHnrgER0mLvWv9znRjlOfg51
Y52zGJMjMhhC/znL2O3Y/AK1gIQ09iNcxzsP//9ZAa4JFLlAgSM/qVwUQp5rmGLKcevaWHqJ2GP3
Uz8MiCXrsq6LD5/CyrbcfHFhix58oFXfHvwLOCPPPq7YocyF5UUFOFTT8FMLSu9169rm6N3C7YiR
aIFVUCHdCiyzwH6CASKon+miHB5TPEXH5drmEsu2O66UQpI5Go1ZUR0HYUEN202qlAlGqkRu5vNG
41t88R/m2lQrsfCKhZv7ldliPXpykulU/QIA+jVKeNO11HJ1+fN4IE0Iho2uKhgc6PAss7SfwxWC
K0ivvPkiJZsoggO8i8t5XyHO8Q7mkeW+lKd6I/x/ShRUzSbRm176WGTCiQuvh26pwqrQqkzIUM+G
K8KuMW1S60Y8NETZC8K6mDiuS1hT8C05olVSDqLQ4ctjGJIbxwuDHU7wMBnKp5VTi26owFmrhm8d
KQ6ZkyAYtYwN93YM37b1EyVX/OiDnC+k8v6v1a6mGV9e6O825/Y+NnqY/SBU2mlHZxRUMBAxd6xG
3dRA8AAdFqpAFH4yDIe0GGTE6vJ0DOOBYC+FcHpNBqX6LdeOUFWh53P9LDOcZ4qEzSrfjZQP0L3T
CvPBdIz1SWqEE0j0viHfFtsuUNCc5RVi9njLboqszymJb+M3svGx2eV89BrLVX+k3Qrh472L5qET
seGMERj+a8JDth+hQdXiUohS92OR47eldbdB18LYanovEXxguaTdUOth0bNhIGHz/yktPDdTHCfQ
qpl3zAL3/yw10eLmyE1geKqx20MovuihBZz5o0LTR8C3TEBvxTMUJp646SEAROMQz6A0+ioMshiA
qjSFhgGqpcrbRm7LGta2FVXzZ1F7Sn7J3C0Ri4LQ+yB3v9VDJCcwmJRECjXqnlEkA+5WGGl8O9TS
dcNONSsPSJQ4e52bqczL07CccQZQZibvzgI0JrJBLVAnfVXNaAhVW9RtVl2Sod3c0BV0ekg57nKp
3dPSPt07njdyWsaE0gFJifgwgGeDvJs69KLGc7S7hFyziwFF6Fqtyi/SIA2NAmq/187uq4BN7xWL
Bw+PQXIsllaDZaun5tJYgSn5Kb3/quS97GZlXQQMgYYCD6qNnn4ltCYFfjSLxBbZihgfhwP+ndWv
V6ba1Ckfck7quZBdrrJFny4LKu3EEgL18HBFlFsCkXmsGSd6alIkah4manQ7y+qye3IsrBa13YUe
Cm630ppq9M4H8azSJEMbLVtGMIPLZYeq5XMvFo6+vESG0NpqwrdtXiFQgesA6LYRkRDhy/SCPtXc
UN7WjyboTTXh9A1jzjpHuOyWhtjgq6KlLh9Os94hZAARbQ5xydtt92W3vboMDOgO3v7/8v3Ixldy
8Q42ktkikozCXWsIjPSlQu+OTSh4FhmUwX4B95fjIINf7p8IQCpg1QWFeVNuYj68/Uyzkk5VpgbL
3/AmoYl+K4DubaRjxvFdu7PQHy3f3vfvdQuA+7CwC4Qb4/lqpk+WFAX5tXI2TsW2IzT5EOErvM6u
8+hH1GmXn1gG5WSOoiOgz57xhybIePQ+B11lCLJehp0ajH2D0HQO6PMR9PtzCXMXzVSW/oNioM0j
yu1HgMF5wKbd8/uib9z2NB4R81Ygr6N1LOJNpKEtAmvU3ewn2+79ErIY1WvzgJG0fbai4RXPT474
TnYf4sbRRUamwcc4WQhHtjZPDTZSkeKqxO7j1mKM+zQB0y4nIspMrpQ440QXZwBQYXJAgplSB8yY
JCAbt3jO8aEVADri/leXg8c+BOXEjIZO/cpXKaHvbVhCBesDbuxfRlZOZbGeqxsqkXGpeYskRxKT
Tn4i/2z7x2tzrZWu7Y8GvO1jEWLP6BC4GwAP/RnABXvUmSahxo8v/LJ+rj+EyDnMDVJgZUhzCgiT
2CmU3wHRnWsrOOg3KNAh9RQVmfQMP4SkZFd1x3CtxflNVumuCqlg+aaKteq37+zRoAWfUDfLad4N
A7+ojYrxp6KqRnXkps64cbqMImDPfqzgBIms/W1cwI7L0PKoiJwYmFJNseDqhGg7aHjgobSVkibg
tiyRMRMD7kEBrGgF944hx8c4D5z/dCVOvxdQ1gebN0IoXDBYf4VZ2TWLUYwCwA7kdqpJJUcqiYpK
twV6myHZ4gGXOlM18A++/hH8OoNbhsrVtLuy4MOfJdeHM/pSE3Jx0XXDNxE3YggpQvVpUAMf4b8k
pj3yHapJ3JF1kRqQz6wL8hvEk7i1Ukp/U0gzJnnvxKyl3sQpUua8KrM88kIwPcA+ajsh14gbPjOt
8RCaF6iQaqwHCNYkA7anizgZxwySt4kg/I1vQZrWPNUhJZJamuRJRtW/SBsHjW3IchSWtnDIj9Fj
JTV2/XLE9WnQvNdSngzGX85GVk3hl+iDQ+Rxzhvk3FRJkDUDlGIa98dTwTvYxiPfPsjcHeCNtSzu
vddQIws0Tscd4BOPNppKutDUheVZok5Dlsz9tK/XD8LMKlmes1Xum+3XaRXAwtvRKlro8Tsvhy5H
1B1ZNFC9mZ24ziPNy5Y2DN4KaIz93oceH2pcU1TzTl3ADXr1NZa4sGOczXHtueg0YOjkkqxbaBj8
zMSU+4WeUQNF36GHpyAhptPsx6s9JXm2uKHSEyTB0lSzsyUyv8m8J3aDvBdwGuZJuHMthWVDhd5F
mWVhhoOdTlc0fvVfc7imiEnNq+B/TjDdcD+/o5IoXoDFslsCE3wPwoAZ+TLbTOTN6CLNwxspV8CW
eC+jE+gff6imNZElH9e8kXlfviLvexmRo6DYhiiV1WE6d/FcYJHNHnTFcHdkd/Qf8TVv2e5k5Ck1
esK0ZCzleFM/9bfkeB9GVwcb1Whjje4KaN3fisKUXAhwOFj97cRYps/rI4DRtg5Oe/Vkc//DZTxJ
0gQn0X7muvanuBNSkgmVD65OBqnI6lKoMSFcuNi8pFeLGsfVDY8eqr+bZDZQanIltcS7Z8+sKZBi
8c4gtgnUNM1+LYzDg19aZfKUYtuub1rFDM0RkC7R6EqO9lXyAw+u5nawdvqnFPeHoemW3LtH2fzR
d/Iq68yuK11NmDqJ9fKvRercfDSVSjGtq+EsKgQWVu411Ucl8//ZEOrOY8cIgxZU5jIhwSnhXCS6
gwtA7mjY2g9rDkHE8w4UG9FTLQO8W/49ELluEEL6khacJgDxtWaCrfas1nuTNBsTugYY/5BHGupe
7VY2BC9Bp8Y56LBNz9dyONbqcVnoX2NUGBnYiKIpAnWgErxJ8wqyzj9d8LCB6haDR4jrFnIMGsRu
dUntToWReeQ0gvsjjFPcIFr4gETGlIqd9GFW0BeuIGGnb3GpAVdHm2CAXTYLK81vzMQtbMfCzWxD
4bC1ZojdoltT2u6/7yqX+BTDNFjocBIWAtCdr16Ykhu+3xsBAaFH3Dq1GJQ5moiRcVnPtP2l1Ksb
gtEWWPVlgNvTtidfQAka7ZqKIjTEyMofk4OAuZxsXniVumuz1XmwmHuxybaM5PysiNP5qOJJBj2g
TB++bOKL8yHtxTKWbFUmNBnUFQUATIvBXRffOuMWPdvyn8e8u4j57mtGCnHHd0HTWM2wnptdByxn
GVqa8/l+QntlYRAxUFUjbRQPxMhPoPR0AfHVL5H9s5E1UJ5TOclRly0IWex6tJbK8LQaRLejx+7t
JR7pZVvNL9qI1T3AjeUwXNCdwP9f+hf2372lVqDFrlyOikFnKslEpN9BL+U0OPAe30UFbj3e7VJe
PsBjQxbc9T3PaOg4/Xb+1uRJZry/QMJC+VafCIjCpXballmIM2YQiaTilQs7nY5DCFjetAtUyJKe
3c84Wl5es84RL9fEmsTbDJEuELqRZTAChLTNfjmCLbSQg7T6N24c+C8IOll3KtuppwoSX7x4xL+j
vVWXi/v6VDDvLK/LNMnJBQJm00lJQeYF3SwTyRKsl1LCrG4v8Ji9i8O5niKnOGtJvdnxj0odAJxU
PMae2GfrfN64pbVOlB+iaXoJBlVRxq7XzWq4h62oTua/XnrHbHZwfx4fG2nx30OALp+k+pV5R5Lw
8VA3fUesq1PrF/4sx2xBaRaWY8NcPdB3avW043UB/xCQpEQzez34Jrd73cW1PpRLNFN8f1dbGPxW
xnXTZ+6iXTKZ5B76uloqopnp/kO/ZJswyf6vm4G5ajQNq991moD/HyOkUYBMq5vSLoWvy8gs5gzJ
GJ50nxQTVH+YEKbwguuUYQRJaw9/2gV050RUfQ4nZBUSPWmlFATe3ZYQCegk7d2T1UdejiMUN+Qe
gGhr2IuFvA9SD7PGXR+4qVYYJo+t9x/pICkWMgiR1gI0KrOuw+Qbayhp4QVLmKbwim22g+dGkKD/
Mm+1SdZ2DXOFbZnaTGNeX8Y4nTd1yyC6hefGgQQTJUrWTug6jbyERussQvhqwJtSbu8BGuSbbELt
wtPRGBlIpu2jGlp/TQJP5gQlyL+B9KKSHOSZFjkT4qUhU4QTcjjaxNmKxkukt2ABkEQ4q7RD3rWF
AjhDDaWeNFNJRMdZR5o1eWD5LUPlIBkw+MeUw3f7ukVeoeldBIfxCDD750s8r65/TkRFp3eeLuWb
/rD2i0YLOdGqXlfD+MjAdjC0Z5N8cTMM4dUsvU5Mk9Z3qYTfsEyyVvluICcxr7jXYkPDs6gx+rh6
3treNdGLgudQ1O7ghHuZUgBS824s2LSf8RT5C9+n93E58IfZa2c0KHNxzBWAD8EX0tS9socGSj5t
upuGRn+DX7BquS/VtR6Iz3EUpEpJWibqVxfx1t3fb9+IHwwAcfwCi8pv9WtpPpzwqbliiqdokMO8
AYmEauOZRaxJLfnZ/T6zA8XgBrxWHRNfnChPBjDkCfGv5CvJNS1MRlVQXNSRbTIWHhaVXjeza4yP
0Z7Hoeq5y/c/U5PUtQgqBBIKP3b7pniZ8Rx7qznX82NiSwbciuswfWr4E5RJvPFmSDMYmrAEE0ju
SsoWrEQroC0GkLRT/gAEWI44uzXpmtdCJT6EscEnHHhvMsQUmamu+kuFo5keWMHF8M8wLFb9vdvR
aL03615e9q+s6wg5I257yBsW88Tv5MN0NDNwXBbelhoaABao9tIy1eO0KSsHOUi7WygKmjazPUpP
msUCq2o2G/ypngPyHGjoTU5ayR9OEzkiC3jKh/D+G5LgSAHGU8kTkHDfde0RyJLiDvkzQmO7hrd8
zWm5ZJk8v6K2cYxrgQc3PJwJNdz4zsXvjq/bugTKnnXAYmx5bGDZEgTbGDemTgUJSiu2GoN/kfCQ
dYHJHZ1NyySC/xVmmpLrIKU2F0vp8JxRg21V+rkqlapX0f8jtstMOHmNluJMRox2jnWb0bHnkkTZ
+sJyzeqIxtgNvEFC0vLf8zgYpE5+PXPOdkf9phnU0hjmKEl2OTlIIU6gpftfwpDa2RtQJIIW2brH
rAL0aRwkEeeEgLRKAsr3jQ66z00kqBbSN8DuoTAnu5UG/QfllrHQA9GKXCzduKBkw2AW4ZOLhXTi
vscw/qud5KsDupyHeXbZNiwFUROsNiGA6jgyKS7WJyFOrIEeI6CobQ7+Z9xLEP9/gQ2dUwAQOlKc
0QAbq4ptAk8DBa+YBWHrq3EIMVwzn1RQhu3Yt9uV6pKupstm/AvsfquNOQBWc3Ui4NYODQs0vTyD
tF5tT2+ikWlIGYBuRdAqNR68/K2z+2udft7M/TrtZirFD6uJtrtuUuFK2LwUdwAKup/m1J2BqRik
NTTYSKfVgKu/tLB4v6JJjsVfoWb5fcvLuT2xsaA+I6+A9iTh8V6d8xAI+ziw0UX7Ubmoi42YkUYX
D+JOn1Kc13IsOtNCEBtxZQRkinRSYdVVz1euqN/6YDIMe4FSrjQXs0puVzrzoqOLuymq4aFwt9fx
AsikGqLz11jf5PEDwoqz3OvFIMgKJwYIPHJNf9sGCFjxZoU/sreepIjRxiq1Si6T4EC3s2Pn7kDU
0ijFQP5qFFXR/L4Hs/NXfiiNI9faa8D1GcFxhPM0dJbOzh4i72zSraCRQAd2egBCeHTITasmbDUT
sXqoxirvRNQJfreYHFbPKtrewv7bB/SzGD4cSlJQbQlY4DmrboEIJ5L40h36JdrclFSZQATickn6
FFFBO9Bh+/rxoKCSkxiba7roe0iXz9WUcX4snQ8SKZzHCwjtU+NhZK/WxALZY2wzWaCmm9KINX60
3xkg32BIFoo8NUN2/2mnA2OdSI/DOTmuOxfSJts0aTSfk5RLhttvUG9Hff5gf0JG0/UIh+KONtSb
u3J5z26GOBP0pdsptVlHf9M9u/3TyuAbLfsQcmdoOVjPh8oMrtzrMdo3EiZUVN1PNGbZ+9LEaKmS
WMaOyvEs+dcAy04O/azXQ5B28bGMd6IQspFzXThWBV3sefLDXofCb1QsZfEl4ajQ4UeZ65saVesH
Bi13B6erS4E1bwvaIBX5+5SUyDcgQDGppS0t6c12dEihtQztx/0aHMGvLZkl2h8zlvxZ7pxtF8lL
a+BZvgKNydescbj9x6wvD0z/Uqf9EcIMYfWkrBNFLLa3tvd//vub2PTnrWJ6YJxjUAM+ZBIbG91F
+RVkOvHhEM6rMT590SQm10Lk0MC7XNuA7TL8iBiUxAREJJ+/YXhgrrJ/1HZWNa931a1u/44OCwfY
IbrnnXPmh1I4aHxHDEBj1K+TtZcoXlqPZ8+GV1FJfeKhO0Mqj0KvxcXH0cQrrGMBX217zsKuFWl9
0+TMezRpkWG5zsd30rWMONo0IhUIVk4qv2J6yAPP83zBPhkfF654f22jrerdI7hB0liQNNh/B2Xw
o2qBAFBoCVi3I+R8NA7O/CUtSZAfeZu2tKTfN2TXwXffoj5Pf2EGz3v6XSRrGmMVySBptuL2VQag
exLdtzBQwGYI01wktLnUdiuLoVIL02lH2KpCSwhNGLyB8vTLrIiJIvIc9am0jHLPJIrb6GGSa/ox
HlWY6/OXPVlNQ/osWannphynnQkkAWVMamCbahi18XLfSBuSlcrLeQ13jV+Htdg7GQ5hhvmpRTJr
o4trxW9R6UpCHeaduRLsUO4JqBs05IUIO6veq+/g57L8zDr23m84gWZ9Wog0dtUjYc/l6Kr0lP99
zMk9rNGq93sjD9NaVCs1EmUIQlow3vxXtU0gXjk3fFeCtNfOlZJ2IJshDof1x/4ODj7AscaurVsQ
eyL8rCqKe2a4GgngkFC/qIELCsqoWiAZvI1rCKb5rJKTRmepWSTdECq/hQ7u1OAyp6j/e62s0DZU
OlHpBaXLigSO5dIWXg4Ds7MXej/1qIktagsav8qbtbK2mL3xZbird91q38ygPqQFhmTFKM3DLw3Y
jTTF9MIwdWLLni3/h88EmP7MHHgkgiJWFqDd6nVQEdkB6sMdQ8aiZByOz29z/Ncz10ieH0m+eZXQ
ZCPsmcdE79fkY0Bg27PknAVxAchHrOrG2/o5hs6e8gM94djCqxRJyW/X1TttTLqX/nZLKZyspF3i
ablQ9BCX1HMms+/cwjU0PH6PR+b6Vhuc7d5xfP2tEPK93QHV6sFBhKyN02pdINHPD2ItaIHRE+ZW
s1lh/9gpZI5tjQ5sSSQtNutbx6C18tgsG1ZdS5akC7joEuuuKBXMGM8n6O6UQCU/U3hiva6lUWSv
StLBHCWQ+hZwQUVuJkzot/1syT4/svcea/ECY+8KYJlrJdtpqM1bb2LeonZbrY8hfdoZWZd98TzF
hq4buU6eWzUOJs+ILK/i4OlKUpkytX6pP+HpdMESZTv+DcKniEoYjT4EFiSYna1W0JBDOI02DCqK
Ax19p34kl9kNjwiI2vz+vgTnTpCt6DLs3+6X74Efo7jFYb1/Y7zhaxc9CXwJEBhToyP4vyrDB9kj
uOQWBnhkdFoeUpafU7bQyH3BzZVOol4KtpWkPv7QL8J0ep9sOfb0ZQh+KRjL6Acl8780u06LChi/
bfQMycI9yb7v+kZNowen8EfjCWPOgWYOlRQ3zj0pwkeYfWmR6XK6LBIzEYKnV5v/jsdSEHytZPcH
vRCUbr+vN3vLEVSHlM1Ma7UNysmeLC+qkM+yLJOlrbRQ5vTvQCLqU7xnk7RipAJAsy1r74oQLUVK
BpcDbgbMXqXvEKtGu6F9dSLvYX8wVkcrVqa/7w3EgwQYbEzrcX2kCgQ0SueiRG0wQbasA5Td9YcC
LaDDvlXhdiqKLjpqS80i6o16GIyTkYLWTFQmyfVDzltDbVuauM5bS3ZXJ3m7frmArcqGr/TO875s
wDuhDHri4+M1/XHQlV5CPIPZknFx4uMjEwmBWZTbKvJxpGwzGOYiOAMKoOQDUq6mnZajDw7j3cSV
VxnEpyYzcy6zdQa+sLtzx7wBtQnvCAV6Be3HjBQVUTOAj7Q3kfdYy99ddaqREeMiYNR/mmCzhxlG
0hco05cR3LbAvUwmUE03q7rIkO/4EBuEEdvmodA595af9lIdyCECI24nD4DeMURJhqdtGmNoMVOL
lfkkDsjEjzFy390KWVYOULHJJXGTm9bJVsUwjVWQHrEtnIn+F6xcYOi9IhozLFFwsXoDjuVFDy1l
nXRZ4pt3dHmeFYlvEuwf9oXC2h31lwXx+8ICLLnLOmIrxgfT/dCAcMMq27FGxQhnqxSB7txr3SNt
PPvbnZKo+W8YEbVleEDG7gB4+yG/kkYwgJWLKlxMtN492Mw0v2LHwpLn80j3zBPZANK1FcLjeo/7
4JQ/Wa8F9IhwyJ5Z+YIOtQT/9TjQUHEtSiaspWD9ZM/zWpuUmp3dbfiJL00yzSkcP/HGNzSYJ7DB
JxszbKwrrH4nnR8JiqUTjZ3r92DQRgUkzSNLZWu4GknujqYLAyyYks0Zp4w6AduqL+mNHh+6R21p
N5rmfrnlxkLwRbMusiLfBXTxlwA4JAdtF1FzPhQy1wMvV8tWNZxLHubyEivgTwO3+wOGol1jwYt9
j162cHMSSAiyEioIMDgLH5Zm85POhBWjJuw9O1FYBfgw+ewolHTpCnglTCX+39Ngazq75RddG478
Xez66ar0Y9Uv8oK6aaGqQr8O+43bNJVk27WKDKS5tDXTm6B2GTWYUUsfQMKNFgTvGC7Mh9+9VR0A
N81ZV/Z5EvcGh6ayxszTwaDSxTCzgPlQMyc7wvw3s0daPb5MBMuFoKEAqdWgdUgg5kfOHDpNCsc3
r1EbuK/wzFukIBtYTLCGKXSoXfGJ4eJnp5LhyRxNShWML0ztP4C3BPDJo1XzetaT5vn1z7T7P7GQ
PELbUEzDQMLv2diznrdASkAoMKemsx7BycpQ8vmganevaFuosx6EgNXYITEv/RzB3r6HJ/J70SXy
stH5iGyKXo0Hk0qowyNwhMOzG73GNndOoSSDQYyRUP/ruA4OBnWJUNeBAaiTLCkDS1hLasbYU8ms
CQX94XLHJgGQJ6pqq7SrA7RD26AYxTFj0F66eWgZ4UN5Zc8Xd5Fb52DJ2lbXlXSD01nGP/Nwi/tx
Fcuq0JwJ4qajQNHaIg0hjgjKPjVaMzgLtV6Kof+ssordvttO9YtlFBJLTRoecwaDRbYGLvB43OdP
FBzOVDdakyXDYm4/gg+IXGMjtA7QxU4iipUZ1fIf8+l+qS+AZ00fiUu9xsnTc5pJdOZ5nyAT+L4r
VT4U6bJ7sDiO9u+QnX2fZw+uYMCcv3oSvniPWfvSa1Y/DBGjnc5gY1NFjYZDgMlP5XZXFvoquDCw
UzYE4UrtCWAcjHdVZDfXNY56GpjfHq9Iwo+8Pze72VJyi36ZUMBGz2Qn+Nxwh3DpzXfhqc6uiusq
2e/GZuOzDxfiB9V9hbKwzYRDJ23p/KVCPMCtKVEL0FZ47PWFqUT48YJtuPkXsLrOnc6q+eifcjvd
CS6mRZDRRNYsOmuKEpw+HYGxkk5Sl9DUvCBMFxh6KzQXV80PD+yqW+KtXVW5OHdt+lLmPs9my2zb
2KwMB7EvoPFzYIApW8i7TUdFmJlp3WB449Gr0queuRdWHy7RwZj7+FFp0qS+G4IdR77dtvHOtwXV
ZvoITmbprN0gUjh/ouSoybIuF249qK6mc5WKPbbAUTuOQaEFPpcmo7RGkQh1/q4ouhzBgm/bFtsm
PYsabVTEtcG8L6YcCOqX+AajVZl4aHtfbF0r7Yubpew7eLdNxI1RQTXi6HrFLw2C/w7eeSj3jYxN
DJfxvzPXPEBqZvYB2/sHsirqxpahbgxg1Z7GjrRaI6uv9baAN7QeWD1/4L9qC+WZpHzDPXsACr9J
/ZCk2briEJFgxnqa0NxmnCj9dqLKyiUZxmNV5gIuqyDazhIqC2/ojVjfC3ZvsieWt5bzrcZqYg1E
UQ1bxCQ9zjJkEPPmFodcbqjsXCkim7oIK5/RLAW4SQduGKTKSN5HuRt2C3h1Zd1BMGwsGyvrHfhI
xUfgeN8cs3+JAaywSOSSQI80gZGAIOax/XYse26wJ4bTVZphUdtQ15kcBOrVLuAE1SZEKtgB29gN
AAl7w72/rv3mG55RsLWZIoGCvOvoZivuxbCSObnneZ1elgHOg4cynTFcQQD/q5YTZNNrrvKUYaje
0k6h+vF8+Bw/XHw39bUpA7rX9H67EXINri79jJONgI8HonfMVU+CeWLaAwV/QsIpRy1cQN7aCEtz
QOZujfw01Rgn9eID9pxk4tmPP2XWIVmudx+CR7IfE+XpSS7zZ3IRmwxoAHSgil2IsWmyZQFEhRpm
1MmsC71XAkyYrXJ/0Z3vh0kGx6reOf0XGV/DCptiR006vaRbIoe4hrLZgGHGG2HJqUyhdOfFSFG/
2hpzHORfMoVG+Z/zyrIdFmquD1FRPMHAo5m5K8YYWQ3hHU1vMY9N53CaAswJEtAv6HlGEMvZrTcu
h2YiXjiygC1IxG+pswleuSA7IELTriel3iYuZ88ZULerUbbn8G6EtkVm56R0n8x3B+E66bJO9WVL
GxQ+L35QumlYf0A3DkYXbxaAGoWbrgx9X2JGPOYr/SzKaXuRufnIqqwlM71tpXO8s/r4dsTs+pM0
TWU+Z6bObU/kMYsPngxEWJTxj/vPjC+mfVtCPq4fluMfHvUi9TkIWRJG4pGnqHkQBTTOz/pfuYJM
vT4djCBxPeqTBqhSa/rpp9C9P9IxKGcJu9QpXU9qK3MZjxU0ekG8DmjbUIIRiUlPEVl5c5tXRmWE
IbWvUmfTpeX2hICviTswbPeveDc2LP1SlI2ZGn593n4qwKMrv3bTVVolYgqKApeRUgFSNUPHg/m+
ApjNzzGoH7acW/5tMxc1gKtCuSxkpPkaKrUTqDhYfWBWvyucXzA4pIzKWasyzUVHpPw1YqR7Z4o/
SXpf/JIzOm99dgZmRaK3LPDldQ1sPVLlBQK3rOhv8yFOGrpl98cDQAgJsSmA02xRT4riu/y6YBEd
vFSG3a1/EXC1gAI0mLV2syZ7jDZRvizJbZJnXE2IV2Yt2D6M+b4JR/x+zRMQz29SLOuSiW3/Fwe6
fEpH75jlnU44B/WR2rqvRfrTYvVC1w2tQ68RZBadglKwUaeIXwstxryGbK6ZbtBEuRRBWZT7nkXg
dzKuJO/ySWMDCYkguWv5SOJindWGKkD0qmlRDqEzgeWm36ZC9T3Lt+yXBBQIT/DddZ995FSdnjZw
EILlRc4t+CcvioIsY69/HSjeydvcx422KDYptF67zv5Wk/0wA788FTbKMTmbc+Tq7qdGZTEmFjUR
3jcAIm8A05mYxptTTboR3PdIhYdcxQMjICojIU++A1H/eTH0pDPozy3jCvXqYdFsnI8goBSg2367
rRJh9ssbolRrMw2jnz0G6qYEzS0VOW4ApgFWWtmsLSd6YotqDntX3LMajRyln1l/1b8iWYw5o9Op
i7l59BEb/aauIm+O1TjJ5JeFXPTI3bp9yw4NWtScOXXKwWs1H5IYVhpcs6naGjIjMiEyls9ogOY8
1xwHombuJrL93fcmmsRyQFevvG/5mpNMX9qUcIqdb+lkW02BKPLCU5S5Uiv0stUPCvYCDPzHgy6Q
bZGXBnxFdgZ16Wx70+nZ5hjdPyn3burOn5vUjqxvxnSLUVqwt3RkRHxdzzTZXmwNrt19HT95g1id
/1ykqlONhlEWNwf+X5LT67eLkyiD23Vo8Gf2+vpbYNEAWiSv/NE5YSMlmSCCjPPDQreTqQsXRqaZ
vGyn3MsEPO4cxhjYcyFsrl++FNi916/cKYz/SEsuixOcCEle/UIoOjrAUhQH4oYCXF8w/xo4BAtZ
1yYcIHl2GvofMDRz+UTE+T7u7zNLv2nT40t+bB1h6/V7tRwQQJzWgPUWaMSR1tCBRfzWSvNuyZBZ
AR/MHfHjCWrtSmCqCHq2ciX2eFXeD6qlySejRRjWJdSNG7De3nz+YGJnmAS0ehFwECOo8K5pM89P
Ls9oZ2KFjlUOqpjPFMUf9DCWipNc7o+J+Srf7psW7G8jQnNBIkyy/lHZPe1n5m0R+542C/aPqiwp
m+JE9AeWOB2+hfdO7mq8Zd4WWN7b65K62B3uDpyP04C2MNx1/fedFUqHpHb8uvNs5GA+DvnzA6h6
xEdrwEjxDSG/OA/mqDxHFxWFBMp0kIhkbiDztO/2VUpeAdf1ydXyQTKmML2UGTQiYrXkF+YiLGq5
bua/HY8GQLnCtBHo7CRDZDcotfPmjpgpgudDEyyGPOaS9U6jAl9dXvI6BRL3rb5mqxPN0x+HHvV5
WnkHTFtKzMaqDM9oj4IDJlR6d9unrc2So66f5c7tUizVhWGBsB8PUKq3h8V1LHDx5VlFjQz9UYwn
hNZhV24RDzBwa+jSAsbqAoUE2IWDLQlwNto3La47adTEMPhRcKaiaUdyIVr9Dun18YzG3trBuL4u
ZB7IZt97QhSK/cYJBvHRzz6xT7uubWnr/VvxY2eRPEMwwkRkelhbIVbQtcDTc1WuiiqDV2c+CsMp
kobaWgkIiRefvUVRno14zOPbWu4eF3tKr24s8WDSSKZWyNFzwpdTZD3cf/kpxEkOQnEeYE7JhyJz
GOic8fKWC8CeMSc6qgP7LZoRS86Wav1jBt5U4MiRUwN4LXRTSM6sZ+Ao3j1HEFhqhvdwJv9GWmLU
ZL5+ExFGRDklqYsJ0hl2aopNjxgLZlshgcgfzyTbEq0KbHGBRJrbvbDeV8JoRFFKCTWETV27ZLqN
B6yyhnHHeuWpb7mdJUmp7/fgf9d5nwUJM2jKYd6oCLZP0SAIrUgy2q9VY7G/8MEoMb8HagVtjMqk
ee7qZQlGssoAbxZfldD+gLTe5klFxTjC6W6rN7b7KojbsYH2VyvfTaK3QJ2HObHAIN4M3wvFFKv7
Z9wO17AkiMIDz0+406JJpa/HQfvMs+g2QWa2GTd5Y8Lqp6Nuq0PvwXhUUFBYEqD+TSnP1+Y3UPgA
glpRWtjVp6Go4jaW3V5OIWxAL62PoLSF58W0kxVYNrwqoZnfpo+fzyVp4bUKrrU9TlKtwb3Nv3jp
Z6prHmfAqdnrrAvBUhwYl6znO2wUV64DPENC/0YpRj2ggH1711jSRCS/noo9EqR0akOy4d6tnyvK
+xp046u1uQQ7luYAZJFl5e9yOonaBx9YHaeE4czDNm0GzhtrSKSYx9fGQb9tD/xZ1LkBnc1hXdYq
mUHOWZbL6vFqUSGK1jOZzbR0iBydXXMmXW1nUUUW84AoNMZPEgiP6SjnzZX31w7F0eqHd5GmNBXI
6NJ4mrU+QfWLKWf0JvUB6dtkmsGiYnubD+DuJOB0ptDYvwAusOLLpYyYcWbVQiWAj3wf0YseByrI
xfpg49laslsLTy9K8FELyK0xDRk0/Mx2e5Czl5gzw7IzyNjGLMgQmzc+poGP8EhLSMhbSkycMkSy
Fri2BKoHlQyybCz0sImLRjamRgkyq95sjQRm5WZdgSEbaKn1Tavs+rygCqLp4bUj7mAUgK2+5/u4
QAb78CH/n6Xjhs02nBUGiWBNlgKTJ6R7VGQMSWuBuAwFx93s1iiE7QCcDsVGMEVu8AmHnh7PchyC
iw/Kq2NI9kj3CN4gF6Ck+BuZ39lxsgu4tzgkgIVCgAPE4muje+I6Coi58dNZDJinLAdCMkuWHZSP
LEhUmTGr/KH/LbYWNRy/Sh/p6aoM6p4djqTcGQhoy01t171hvERumDBUmTqCk8v1Dx51dZAPjHDY
G9cKWCUQtciG/tgN+BCaqffJ6OugUoeR/VJo4XgoUpsQGNiinjB0wBqBvo/SvS6OvQ/b8HqKr9Uh
GGUgZIqNThuwkyBscweqqH9rw7C5toCZ/Rp68444SoxnH1AB67rYFGeB7Dse48czId5Syz55XrKJ
PxCiPallFfI89r+ekRwA6yyyMQCR0aIX1CzrftySbcjQrVgaCA2jNOo+2bCzFqxnIZPiJF+5kqK9
R+0DjDDfJg+TVZSaTDsCJL4tOPOyoIYYiFSmPdZl+Z72CHJs6GRgzN8Zkb6riDMffOrivgknaRkC
hYIVdyrzI6Vcik/e8FVeHhJXVSlg4yIi6fAQbUBxSbSQZBOkl9LeSyFu9LE7+DK5bfX1jnc3qnCc
ra+mmz/aFoD+wnvrSWp25vnIzmVZWGFGEulhrPeWi0qTtDr5+bGLcyXqo8MB6MbbhGO9ZxFMagkW
nA8OVe3/uGYfUk8kx6xW7QS6aq/bgzs+mCAZ/vMsFOo1JaAeJNQW9eQvO3QKcjv6xUwR6WqgEQwz
Gwk8ktBH/q5+wxh8wviV3PdbppEDsEJmffndIm3HazUNRTVYUSOboFwxURLrpaSfijQ5Ca0oNr4n
8V5l3OA9f13HmupmCv3NHFvPh03iNcUGz7atspIeozDEq3r/RYgRyxMZqtEJ7cHvOSj6VCfKycyl
sQU9R9Uu1oKW0PF1xxwd7FIDeb/zpNww4f+VbFtCx6A0v5Q7I1kzh8iMS7EuJJH39XLiOenz/LXA
0iEdwcaChiXJfKlg7tJ9o/zADNml26oaCzavImXk9RfsRP7qjwb7ymhYC0ojVbZ5+YJ1ibB/teVp
akcfSXSBbJywFApVPB+IAxqmer9oTNBJd3cZCSXT8ucCcsT2G/uYfyjsUKIlKWdxjYxqXsUktrGn
MMr9Mm1scqrY5uQ9k6f1lGg6MwljS+Vdc6nZeVNbzVOIgcFoYmhWeMyYKzToEv/ultzo7I1G2+Ha
j8zI3t1K0zz6PSHJKheAGY4sX/VEueT9MRFhMOh7qGY9RWIW3wUAqngD07WMo6LNWeOZYnciBj1S
Deng5eQOpMzlgR4sPQkC8Pjnaw7paQ28aRQqwinZjiBxcylHRg0JcsjJE3EnnNE+07cbRiFzSGH+
Ug7wzbgVJNpZl3nUF0DzEhicSMaxryNA/UCltsqs3BU4eRdtasJzDzSfIW9QpbpTorzV9+WwuXa9
JpUSttG8a8ER7ug7K7wYdkS6uWFp2cgatlguWZu4nWlk5bltOYJ6kIVY/5ej00FEsb/wbau/gMGk
qAcZ420UeijUXHrKJptZqc38MRYMCsPG7qvCqm1f+yJNRked2A5PxLtZMUgFv13WiV//eL9Stxy1
NA13vsV+qf1IhpuUIFzP3BlB7mPAt+ujNZkgnUz4S6pjeiWcSp2UIwSUoyTg7oNAilmvvQbWFVUw
GnIFVVf5etOOW4x50d1xd9DwuWBbO7M0DOiVVCkp5oI7JkgAmd0Z6jxLKIWVZ3KN0XgGX0AcTuWu
SS+FGUrVkrCJcfGID6bJzw2HtIWmXEqNaYoV2lvEuaakzDAL1qGft7L/Mf6GkHuLxWXJ42q6mxbc
NjwmcVOv+xJc9rqFWPPbSbEkVfvS5WMOmFd94YoEuDWegbykNncx10Us/GCSvpW3Fx2KNcQ+EsdC
rvPLIdKPBG0D3r5yzabBnXShdmCKFyphK85gD1h0knumUYiOjUIg4DnXnI8PXFpiNWnmSNN7dN1I
YmINBNOn4Cn1u8GoreT5mjyrx7KNTp7EbCMXAWgt6ra+lTnwheIeI/3o0ZnKcR9OgbTQ5aD/m1G0
fiSSdVIL0giq1Eco0xCUmJtjO52dx2IJHCFLaFqJWx+IAzDXqwqdjkmmEAiE0lweSLSUvftXnwlL
LufvGm7Vl37NzgDdIDto98xyDdpOgxVDY3DYSe5GkiNZiLpEsS573/C2zn9x3zRN2zGw2We+LsWV
I+Pu0kdvvBIYrbQF7MWoD4toDpUOcBqU65Ef/vPhPfLO2C7kz3AjBcFP7pCY5VTXA5u94qxZRsk8
jLg9UCi7eei2sla/A1j90GI4GMz/6pYeU/q6UPWEMZdyEg/Xxce4yV58lrqJJHanf0LYgoUgQQWb
4CrMcukERLT+TBQp9ZOVtLSNbiZ0Xp+c76ADODpxkJQn5Q/HksQjephI5XWxNm5SNf/f1wABORAM
dwy3Ildf4EelHSI+H8ZTcfba3HpO5anDUJejEsEruLNRg3dxhlJI4JdXdm7/8C8cuxljinzke6Bg
YPOqvntEPxoPaol1IXYuyJV/5Q7JHLgjcbOpunoDxRs3gh5+m93PBqWns7FtlDdvAoTjJCHqaWCM
8rReHosUT19HUI+W8y9hMyDyg1bmxHniHlP5j6SbnJASHRQULUGCtLenZLKYQLtil3hSEQwHDGVF
U+o1MpknbK8IbPziZRALQMO+C5eoliTKvR8BUzsuZk4+jzk06f+NcCbzbFnI4T4ZFhBMbVEvLVvi
cGW780mF1UvWO1tPHw8QqfVDKxWBy4i3uKtjR9qcG2jLcfUxoYXuQ1ToJo05WvAxLhHI2RqLymlr
V06KScUmL0hWMiO80ot4w+Smkz9yyNZKgLeZ/sJ/0wOGSDvcEi5Tc0dCEq5A4WDcO8Z15Jh2Q/YB
eOhw1ql1jPld4tHbOefDfIj2C0DgA4tOH6zztfacQJs7XHk1MbZXZI0p9jCAM155KqpjzYeNUDza
JCdESiVD/96JYpMEGJOv0TFv9cmlvW6IsvG1Zgcf8bj6+1QTJcLUTlIBKb62benJUyVY2Qg5YMBf
pDBBRghwGGmJxB3HyyGNgHfTzrmjnmx6NZUSv+CD/Vx12LrIXDlhKJHF9bbI5skPqvHUYXT12EAC
XVwL9R4o1U2EpUeaFU/FcgU9GyJDWfnd5GcpgZqW/2kLnZmexXiKba74SiL8HXuz2V2m3JvqCQTm
yQ204s6RQ4hWvxWEIGpoYjZdcm21SyUo6C+QgCrx6qtCKMTBNPMhOtM+u5wnnfEwSgLFay5bf1sN
B2HGslgWIhwAFdiiwxJv0Lzf1sG4diCAz6tUA91/8OZaV8I5xTczRCsTh3G+LgYhEeofSPnHleEI
DCVZObMp76c7e2AL2CjANoZRqwGDyqILgdmK/5GGUisqJW27VroqdiQtWzsFXyyUNJnBnvItEtWH
du25j1YKDarWdoLs0jdpnU1yyw2QS3TWPICSCSHxiXz//dlCmnG9PkEFllSSLfynN2AOBLgdn6Om
oDC6npgC0w1fQfpp8X8mr2B9oGFNPs3DdZ3cc/XSIPYQmlxgY2vcFnVpdgI6qRpzJowZFulQKk+E
evS6clYVBfk25wyUTLsifAmfdS0ekb1JSORq8B8SQodH/iLb7uzURv/rBG2TPQtPoZTZF/ZL//xB
tU+effrv4b7ouAhQuUK+5etyP+dQusjKf7lNC4+0ozj1GWWHasxq28JnJixO/Vjysr4NxeQeDUlr
XKwJTHV4w78tKQfGznL9fZqlO9vdFySZ8EOSE8WoxNNJtrCMo/qYp34SLMNK9P1lLwvGX13/y/39
fydJmvA/asNtNLlCoJJmrSjY52ZB+OCyB2u7tYcT20YehevahIVoZ7reBiO0o4gVwS2IOYugxD5D
Ug+OvhUgLO70VrcOMrdhObB6C5mbMty2Tg5xbZBwHedpOlkLgg+DkfS2axD4UQoIkMJyg2DnGqqN
/GUSak8NEVxijERC6OAnFeAB5R69JNVOWm4cBeo7hSCb1NwN2iKC7wABd6vYtENtiNbhvRb4RTAt
Hu4J6R8wqCAFYMFmdh7IDqhh/ghPz+/tm/+6ofJn0fOu9J0+mErRVPT4gQzGsz8Tq/jtRQkspvWY
Opg0iimlMpapZEQQPEl/JQXtf9FeYUP1G7IKCLTpVEbpJqY0OTnF8MZgB2A9BrqJ2cfNDgX4s/uJ
/Fbg4e8HxaJb4mAiRkSuQbyDjv3/fMP+SO0RQmBgHz3TA++Kud14aPZu12K5ulwKzp1xazDFUN9I
kSXkY96LjHeGc5kvdZsy7nOPpRmRLPat/7dzmNwABbiHKkKGWkQQoy/NfRg0tNJMJVxemCk3Gc36
0DN7uoHDkA/+ckJyIcLxpWAZwbgnSZyX8LIIEqeLwStwoM1AZA2YCb+0bxd6PoLUw3kEIygCEdUk
Mcjnlen1cbrXMxJ1NIMVlE7rr7catcjXEBAaAfu8H43cExUYIhtp5QugdFWtsYaByiUV+Nc7YufZ
Vb3qmBgMPR7kw4aR2G+jcIRjSwHIP0em5MmWX/li1iTSSwqImt7O8c/UEcb0XO19Nkq3A8381HxQ
Y/b1rXowzk12I2PYN5djCgwfcbI1pk9kAp7kkjsoJmQMXDN6hUx9rZx+6kdJoATa7PtWq9BVgjpY
OSj0INI5Fb3V2t0OjnGop5JzWfdwAzq6Swynu9j1IiIUmdchYW+PYeu/Ng/gi+U45LktAOEr1AY4
zlwNYdHB+EOOLG4VQQX+rOtTjUPyvUGWEwOWyj+PS0aK3cSblEh0zaGLZmeJzcjrt8IAEeGU/+DS
7wQ+bRqx5JIDP+q2tyZkB417Lpufx8e49DoD7DLFzdX0nYGUF/TF0xcN2RdR694F51shxEl7EzTx
e+LjCtwcIxLE3MRNdXq7PczZ170znefhFmrnVUxdT3PgTbmcbIFH/zw0dU6G8ew+DFiCT7tjX7p6
/pzbPlJczbwLTpxQm6dacLMCy3LVG0Cos6JsbCuHyAN02G9Vw9sCv5zKr7Tv9ek/wYKYwNHjGdin
5ZaCO8fCByEIQd0b0CDTF5yrdO1VTybFmR4qWwENyZhPh88w4Ffaq1HK1XyGmpVJoZ6CZgD7AGpT
i1pkH1vA6QoUMWmNAh9fHrLS1iiS/KzixWemAnGrJpS1ocRHJBZNuQ/H2Yxk+YlrQnPP9UCbldvV
npL41ThWfqMUaHEZvMYHie8GP0OftuPVeD5tq5VNfA7wOBwvaf7IheI4aVPKnYdGFPOglA2Gm5SC
gIf3hO5fm5Asswvzgz8FmMsPBK2zgloWRANa6qrrVE4Xrfbm/muc4F84/BFPbEWXIXWFPQVZ60jU
EWTpCel70xJt4hdf9lNBE0JM7pEuB3XUj8/ULECngsRL5vUryjNlxJNX+87LUOtHEBsc2XrrRWK3
rC4//d+EoswBTn1qB2ZTKDGj8uE4wQlTwKEnZxd6glKjM8Jcbl3uykdHZ6U4BEfCkyOEMFko64Hg
n4UJ4TuVIZX+fu0AP39uXsD194IuGrgzpthrw0DjusoQrJmNPMf/ybG9iH6egt9u/5okm/kz0FEp
eLFaEJjinlYqrxewrwXJ7EBKOfK/sLCn4FeHxO4QDIDW/MuaA604l6jpYLrmYl0fWQ0HtTqJisH4
5ulUqX0RBCVdwZUiEqM86+nrHwAuRws4OXfV2SB+JEunt89yEv/BsFmnuBQkyCO0TNBhDCai2+4n
pWI3XJeottPLVu0DbAtxXiJjkrZ6CjmiBXb/crvEhLmqWeb4g3WTYMWs+jtKdmeCIBkv5I29nYP/
wSMe2qBmHQLwFVXWIJRjc/MdSaCMvs80Zm6ikhjoeta8Wl5q6QnAeZuVwWrxC4foSf7lID1sc2Tk
glW20GEteq6B0JORRpnU7e3wqorfLdyRmP77/XFgCsVQRflmI5UCDWX36d4qWBrfaXPbnA6NjqZT
9mtp+tsSo6UpK9aCnaXbbVddZBPf8enmVWguw91l8JKkEKK9DkKSx4lxc2qdLebAV5CHqOf07UfN
/t6SRQFRNZXm7o0X02DAdtEiM6YG3lJ6SgrYyJ+Xjy/vhVKxf8UiP1o5ALP9szWEQktUmvA2UQRu
9Nt/FC9DA00zUvZj8f+NKqYtkv9lzN5d0UwQ4CsVtzB31GZmnJt4tQkwV592YWg35q2SZX/8mGaT
BGTiypbw7CNLRLjic7ZTm/ZSYEe63uWoOBACLsaWxLgWplyHtiV5RzphHrtcRxNkSnqFqmlRL9yn
2y9QGKRsI8DhOvJWAiKhtjIxviZ1PioBHds72aWsfFKxg6jKbhjoFeo6i25n2sZ8Ka2lvwOnEBTT
jNGiTaXiK/+lpMMh2rH9q+blD5BAysNNxhCD6ezjpmFv/H2WXhmMiYZydVLgTcBOxmHfhJCDm3pQ
AeOIbvfueZPXrmfEfh+pHOPZoQTkzCBX7A4rrbmiAsDRGPhAZo31Fuj2vKxmYjfmxE9tiFKyJk0z
RyJWXfMLBVfboTo5I2GzxXKZGDIhiQwHw5jBcZd+yjmw2bbvBrnJI15S+CVmYqPBYp1c3yYSiuXA
GAJj8Y6SI26fRyg8UoD3gy7ALseij5gHGBlA6qGHbbSm8U4vCSMyBHw8/fQUxsTIIcUD7NlrlBmI
4rD78u86nGKsIT1K4jCG+GJ5MzuKOti9J+0AYHV5t5vrnAP0Z0PepC95lZDPCv2A5GyXUg3Jl6Hk
6YkjkYjvKbLfphKCgJ2dFoa+mFZA1TrHQBUCEZg76JJp9E+myAVcch7fddynwsz/F7MqmUJuc7mR
4LITYQFm6S/mOhqN4WaIUYlydURyH0pZ+iaHRCPwzd7mNx2CX1pQXrbe8JmuIIUTK/G4YlgzcjaU
6g8aaS/uCaO5THzcp2YCy+uqsaTpoB0ZU5U/mm0qj0fWqtXJWR4CZJKcR6fZFf6SWR+u6NGyLRR8
csCOdO1+I4zJrtRccL7f7lqzDtQQEHkPMrP+moldD5f2V58Dc24A/Uni7aREoOd4L5jppoaD87hI
OVRDuqb8jXOt9JHCx3w90T8C0Fc+j/sBZ1+XCCTgWclyqP4XbLA+pPmZK3xM7JYByuU9LVYqf5LE
AD56F7auePxJc37xKWk5I2Gm9fWEhb9GcuqMpA2Kk3wGYNZhYg6lCYQ4SEfWVp6vdXy6UnRZPBlR
1jOI34UAvZEhGsdhZt3xsTexbhvlJZhsSorrRFPqC1/qhHlpCBrm4OBIzgPAbjoSmUtZmxbElAuC
GeNEVnGjEKfqm8l5xgVbaCLXjWAKtdQ71lR4ECecFVIuTnz87Qz+WvtWia+6Wxnbv1eGbyCc6eRT
Lkv/9Tq+RL81hVzrrKnipDC+ubr6Gv1HU/IaeidtKvNFaTTg7J+rJRE907lIuT/ajH2otBDJPT7a
59mwPSJF1PZF1dyu+5xsCmbvwL6678k0A4smPzhes5KDbPAkVrscGmjNpeG/PCw5muUTcuaYzAct
9oEt86godtkv6UKmoqG31jl1VkSLyDUqNGq1PJqRwqZ6pe8qN1A00jiqNADPducyQTyVOE80bw2h
vSRFeS4XDCJmhkb+eFByhqjiWPIntzObA655zkevOCaQzUm6Cd6Fy3H+VWYUUqNC0DcnqVxzsmi8
kF7FE56NXaAHUslFl7wv2dJ/dgbPODy6hWdUy8VX174imdbi0DjuwcbrhmwaduizLWYJ/tldL5mt
CsnSyEifZTsKUUy6FeBgqQ9RhKUrgqWDb38ah07S3fHEnR/RAET0zdZKQ+PkyN4VELzfFK8Em+D0
FsqRJ7qGcYeNqj383aiWctMBDZVuurizFpe8lBKAKljKUV8vyRyapoXZtkNUS11W79b5veWUEYz2
X7wXATf8p7Dl9ZIB3As8bnY1PWZ9gRROPbcg3aNf0Y+YD1Yz+wA7QxRRQrVfHztBHgYg2xtrOYMu
MHiCLzb/fN8WkTg5iz5vlAEqcAjX1+0M3gt1syVNjxE4vFmjBNAluVOK53RXSGNPG5Q6JJFddn1k
SBdboDcI90bGerr9MPbH7Dk9bbjZpmMUVWp8vukpiGnAoOxaL2PE/0KHBrjEXOpJ1kLYFmx3i9KT
Ftrx2ibYf1sgwTu4f9Ow+0xgLkiQk0XiLa53W0gnNit4rKpFYbHX0VxJIV41/7i6iVstCmLYjaOw
DKz+fQyu7iDqMhOtVf3ResalQVmpA6J4+1U3I4sJQR7vFixICcI7Weu187xm2XhN8IzC+utkjatD
/gJMyJgdTR+bO7o5zVG/12Z0lfardUSFXvw9OA2lI8XbX5OqAE/eNnougZuzpxw4CGbnlk1fZ54W
23CEQSrxMflgn6Fss1eH78b4skzx+mtGRszJkYbcs0rleARwAn7M10BnD808iYtcY5TusezpjQaW
xqSRlbP2PeVHwCEWJVj1UNazyKzsacOnesy+h1guJXhdcCPM06f+dYs8YYHZMtyi8t5vbSi6DN6q
jJ+Kul6VGG1BHe4BOjahvkxXQ2YtWrtH7yCxoJmsx2TDAn/LxU3r+25HMFWMUnxv3KtnT/JpIs1N
84w7M8FurqRnR5zU1WI0u53yI0O/g8FusyA8wBScWQHxMcgj8QAOcYOHiidSzRdl2gCb+KvBdKg/
h4ilu5ytdqVkzrZs5W7Bo75iElShuNUKQWZr+NJgkU5kSJRqHh7k1PSbJNAUKGeskN1JrS7dNlMD
T+JRS5TZA4543Zl5gifcteVSD235H/UX32aJZDA6k5YOdD0LZSU9eiSTDYeBIbkX6YRJBlAJRMn2
oY2Vk/RO71vXX7+1zyFXK8vcwdHA3P8qRvKRXv3LbCWSsbHb5ox38zW0BmJX9SOyAf65TLejVd06
ijrnHaQTgk02JfeTu9/8naRNLubca6/RMg282BUNjaEPzalSRiEDubYO7b3EFkeoADLbLaspaI4W
Ux9oiPDrTt2yRyqvPymkmvKC7RjXfRvQgFrYcbjou12hQsC89ouuzZMeMYOWTNNF3nbWl62viyhD
RnD2MR7JipU5eqGfx79kNjmfY9u8bOwgPLYfEuRuSOBnxjMQrRiCaTHnf9RZSMtVh3Nkb1GlxJMx
6Xr5z5VAWzRuMDtS6MoB+2wt5WFWD4d2mxRDBqis1Nk3EzdVeo9ThM2wKiwKXt/SqL2RUr5FvlGl
R/CUKH1RQ18J8Bzg6jVBfvak1qD7mkyw471/Zn5yrtBG2VlbpMI0nanmrMqujcNmgLWMragvHrFr
IhuLmGujRqWCbRdW4by5vhCHaBz2EktMDWw6OwJ+46vwtHW+4bvzK+i2s79uJspnY1PBiTCo6m6B
8/ziO3N8rP1zHIBFZ69LpuhBIMS2fdfoSgHKfVl5MIEOyLk3Ehl4dTeQQJIV6ILT5DlSu1KTsqg7
ikpTEnLTHUkgwfEg//YzR3EZO9UZgEXN7eTkjRKo4gER2Um0fe6DxmpqJFLO1JyvmK6eclrgzZPr
+w0vjlSqIz698mWxMPEJqM7QjX9UQIr9KRfqSjBFkYvQLfve6Q+Ne+fbgCE3X7yfi8YHevA66RWf
dn+RoM81MyfOMsQYXZ0ceO5hDsY96cOwzJhUv+SYYTjz7Y6gSIZT2eHrCbbMRDNygKyguO35tpAr
fsCkG/FxbM90SUsVZKfxA7t0GYWBXyRG0TXr/7K6KzGylv17bOls7/xBnk7XtwFnMwmkaTovqPSh
gtx6YP5S+qrKgM1oK4GwxNNuau9bUwJPoJKRCRrB+DbZ2qq6UbW5GttKb5e0UPOfejIfsfObwgPP
+qeij/4OhyLeLIWCOdLKgBgmrmOdIjxpQJFM7e4eBGQQzrKEM3T4JCY9XOffN0/9M7KolUehKBRH
HAdOB/5ijK3i0eBWKp8HYM2+phxp4G3m9lWoQH26bWiP1exxBHi7smRnMrYsc4sThzRjaNLFFIQu
t2cJ4e+JnwL3AJtwCnVzlxtlqL7Nas6pETpw3zvVgfzNIfQ9t1atb+3gFGzspuzq6TPh0DGu1vu5
ehuYRTDxCWOzYP7cWrhvYoRsQ3F4YyFN5OpYpa+4x944kEf3oH56b2KT8FgaoCI4BGDKWK4yTs0y
Fl7qjLC27sjd2Bj31+yUnwnwJo8eb3egy5rAiiQIAH3ur4t1Tip9zSqKZOwpEdAdV120o6beTDe2
Kr7BfmC72vtmTAQJjesiFNpvDuNq2Svtd3LE7yU7vmxyLVGT0sstLeRTTPFNFXUOOGSsGIl7VA53
xvynd52hszpcNH6RWjzv7ZaU2SGbd+aMc+UB0ySc4+a9n9Nt+ErADYrsvN2DhAjfdhPqR5K82Afy
q8EVWfqyBlqjc2sK5vrNpVytxZbqkDzSY/AD/J49q3k8SsExggdk51cI/BZmx5aXEfLa2+3JETKn
7Fb1LoHVhe6QpD2KUL5EPg1+ZbQGdm5U2P1Z3OXLWOMFHo/iYKQ3mrpP6juUUpuoqfrKq/s/yR//
zaXycvUKDUKkgQsc34A65XncLD3q0Q5jAn3ruABT7mpb2VX6WJCi3rOBA1bxFcTSqO7RZ9FJ4avR
5fuhdBm/atE/lrklfR6gXXN3oCDyALH5TMUqa4hg40YnzfxL9RyU6o0kE/DVt+5y/3cfnTBeiSvz
L95KMVnopKjPsXU9hSLnW28tnTAoHwtxpsnk3YowKcLAw62qFH4qgESYyoas4P9UphgLyE7osao1
2rbz2SW1ruuUOcbon8yOqxcjmvmoVjcxiFnDwmBZb0uVyXoWLdfkHAqvEFGs9reBsmZpDYf4jBcS
lKQQeQN3/5+na4DTzhLrFA9S4ZL9Ed/E+vGr0K/6hLV59wsOC3psGRpesJr9TkFISSjk+GMZsrA3
ZQjqf6Xnq0cIywHM0n0WXm4Cz7yyjQj6Fcmk9SYs/aautiHapU+KBOWABtCNSHhfqsaz0Zgv54SU
Gg5+AGHP4uwuWSkNyCYno2riAziBQxrM29nUd8+KhKwqzeivK53lmtM0qqzp0yr31dCx8X7OByY/
K8ZsgvMygFtURs06JYpf41BvNnp4wtBV9xoLhZA7l2INFO+Gp68LzuIfY2oFdBLUqJtKLEJcU5Pb
sc0FijmHW7fO8gjBruXAiIu7nyjYCWT/BiBSM3IZP7xiAozxAA8CtkWaHxZSDotUgjSlbNVWhljF
Xg6AhddgUugT7sNgjgc92oF7TByeuC0cCaxH3JF4LA972owIPRSQOOBG1LfWF7FXraFVqHML+L+e
VBBWJLH/aagFCF79AVw5hXyNxVV4zd9ITLFlqCEUbAP8v4FHbkUG4MXt+jXo6FLgrkdkOwzFyEky
16j/+KzPbJhYBJB3RZsB6By6qDiT/RISIavg1SjmaRhkFEBdN2foEpEavrn+EaVDFrfHVLtxQlxC
4Qk46Kl5zs21YBRuxKZNSvObqO3kE8jzA0z+Lby+WQmGJM43w9/f+BZFx41UatEblNZjrW1wjz0i
VGpbZax3A0vYd1cAspKs3hSIGy4HEq62s6Xgu0bJOrbwwnwmk7bqntUrVBOMPcJzVXVsgUfMbYco
5Fv7Kd8IggPGjBtokjoJ9hrYLMEM2tQVPRwO2u74/0XCwDv3A+xihhIycCMIZo/3j0m+QG9ihb+i
TVl52h55VaqKQ7OitCaoQp0DaxInHqqTELZYaTVRdjp3muQ5mTX1sDUogAjQqoJvbMZFo6e4D+Ma
J6EQfYQJg4VEAseyLyr8/aD3b2SwNBb8QqmQ2p3lOfWGoUWCu8WKkrOB+zSpZD/Nn4BJ7ZBeUbZF
ANfgUq3eeTdpHc8jGHU0UWWTj91TtnDEP2XYgTFMfJhUb+Kb8Ofks0I1qB29flxzsoASlsJQwl4Z
JclmEvHVd4X/UZyMZdeFtffgoa+0SbTSnhhK1AYLOQJCBwH9yio/FKp9Gi/7WAbNBF2/NHxvQMvj
WLSBWjO7kf9DdYfJPASn6aTSZ+qRzxYuOP4TVf9EOfcDGS117cejx2Exr99oniXl50xapuzNbo/A
Pnf2MJ1WvRsvl0sw54njKsPe+525tWlGoGSOSbzk1pqPBBFF1mULV2G/KYfePpvKM4MQC7HekVAL
e4JQ1ZaY5sy25IU0tqzf0UZnESZmywTFKzZrvJK1djP3iSXarEJ7G+tlDZ9gQCaHOkPF122KzKR5
HFYMZhJlUKlNlBTsXjAtwPzzUycKWL7Yo1IuAzWRZpp/5KXwc0cf/jkmdTehMIiCY2uNeA7i+a1v
AnQDzDNOVXxT+XK2TtMwVwYhJyPAup9hNcE5GA3lV0GPLZT7TxmCYGvb4yKzfxO3GNenjJCVvUwr
JxE8y7z5u+hksNZZU9an2Lvk5wVcj69U139LsJ6VxEHqyHI3/cO5HngUN3qZypcodUB6EhEsA3EI
tClvWcJSLalcfa/P/PXO56KWHDadNcCyDLeAQh26avMwckbOUAx1BFrAdIlpZwRMUT97wYPH3dOf
2dSA5k858BlxMSUZg5kq0QFx5UhFxPJ1irpe9AGY5xJ64XTPTwM0avloq8V6UkNKZR1V8+d2NnUi
BJVJhPpcRX0sE8U5lH+iVKn20qGLaFo/iXZ9ey8WGUVJoihvKT+OE4TR8bZw/RJEKhSeNcKxJVMw
+Rp9fOfZqfQObagR6TMNi/NIITzv1OlAolH2IXDcVtnd31mxZgblLMQDNz52g8fe+2Fu+nRciERG
/gv44vb9LbD4H0gzId0GNFX5u//Nkmo/yNX/+WHc0bM7eWupQIdD5fbPXRnPh4kf34koEbrUQjJZ
Lw05cDLncCejqGibOE8mRWmnE3GZrPzQibhxEy9i+uUZrm+y6OzGjxIlks6Jb3suku2oygVwvzFF
PI7F0YOgGChGmmaVjcjYOSyR+kRXan9+Ppx6oTGer+7U8DSmpLjfmDvqnDgABEhvSLBbHI1Ns7om
MEd9K9ujBiMVoByt6aNp0wGB0fziqNRdb6qpwUz+9gGbvsDY4tOIfKi7+nZ5jdIkEXMnHb/Lhsdh
zdBchoWz4tWnCS8Ua5G5PopcLy7pHHIAuBZsfQOf8lAFy6oTCFDT8QpqDN2vJSkZkdS+faYnOHPc
wK5o5f1hf+jh3NYD6Aaq1Ol3Q4U5tgfka4KcaNGZpYvaAazW2LphPFv6LH3VmzJDNMfeYqyk+Qip
38qsY8l9U6ImBEhLO+t2sC9rMSegvJtTWptKNPL2z4zQ7HEKoZN9BisTukc/hRzf1QM3+XouA4zd
ygokNTZ32A2Kl5rWZdHMkeIJxTT7THliTOg80ijyy9v+5Ve1c63uvXgRugCqaCIwuKmtb0S91D70
tN0xoh81lqP4QAiFNj7BO9yFOmoqX08PSnS7249M6fhinHaZ2Rw9wbcptFNU1lFTwY2n6K7zvF4Q
CtUFKWrbFGGYJNz6kEUQMcslAlpwuO+Edlmltq67GODsAt6zkoQqJGrVYBrwtWCZoYKYCMO+Ng//
KrByblPqq4JVFGol2pytDwgS0f76ZVJIMxJ7ZKQNn0GZgZcYlWNloQLERjcJVB9iDfiqwILddn5w
/3W0yV0qJk9TH3ZbvfOkOsKihF7Ajv8OMDrBbHZCAOMGG1CsZKpqcROC31oDtufb41UwJtVHdg/1
x/+BRiVz1NeASraoDxqXXDoPelPGFQcaN3AcPNoDhAr5h8hBiwqlqVBMuHTcXjf4pYGCjc86QLhh
Pl5tmoM5WC/PTLqiRvql1zP8nCTLULNgNyCJGP4qbMVJv+Pw+afuvlRRdR0Y72KBW8DPIwDFPH/R
bJqc5koNQUdd4HPmsv1+GGHRKhg8/rGlqb1M9/9VE5f/Txqcxe6aHL0nn5NngKD/OxTGMzeUspVm
XlojHts93IB4C6L3zeNrfaRUGoXSq5LwvPfgc2C/hVe7cngtS1WsszmnE+TcHrXwxyA8fqTppOu1
QWj5+MhDVrl4mzJ6ZVcbHsgjqa1KBcztTkZ0yaM/J4kM1/T3KfzrlWTfSguQJDqqbTKdW6IqbAIR
B4g8HKEWL3bupECvHjByUENOcXyyWX0JfYStPjwi0Kmei2zjVH60pEhvZDE118YDyLqUesEsd/mq
h7p3ZPwJM5rZJArB5MG0MKoltfGXT6UoxF5S7Z3cRaJu6rIL4g0uMt5ydwcR4CuqnyzEenxZMduc
aSRf7ZE1RsSCBfmY7hJYfdvUO5Tbd78v8fGZOm/j+xWi/jE2HNck8iMs5jU2a04/ZLSahfT0OHc+
9n87dZ1HlSX4XpaKna3Cpmm0XPBoAWjdBiNJsZ1YLoS7LXK4O/F8P5gK5V9GiHxXwOr8Hh0iTRTy
jtbzfiqQNiL/3cryvJX2MwGWgLIHEfbYbCvVS9Neo1zuFm7/PFiqnpVT18RCscpKKKHLdUYnSG9Q
ypYDSGfVF2RjaSIzz1SGSkMudf5NhKXPyc4w+ekjq6Vs10JpI9WkCN5feCpO3znRQ1dbwBxklWoy
Alt1L/LyCZCJZKx+2Upl2aVnuCmZQzGlP0cFpIghgAgsVotwq8Rf5ai4PiB45zYfDMrvKRoRrTuZ
g3Jqd7hP/db9FArOIB8Q1GMfg0Oq9sqiajXGNF/UPGR0jWT+yHPn0JWjkXaTXoA2cc8F0VjNSbnH
CmNGLv40sk73zbRkTeVrC1e41zNFDKT8CNaZpdlGCFwF6voWPdOptUTSXQfkh6XLloJHsLsZ1Ap+
1hhSB2rTflfgiiI6vy9PqtUpfwA8F5VzwZbg0WP9rkOPcQ9U/NBJvRl8212vLZM/ZpTJp8gNOrC3
X6k/6bPkXq6oOY7R6LO9s4GtCamx6QJfquApHa+vOgHNV4S7X1hnFWKiLp+mFTSpQgX+cuCTAp43
5SzGoxxlwn8DVGXtUqP2Bg795aAqUV7D7DP//qSQJlOftQla++1d977upkhz3b0DpJ7624VGmPam
c6mhcx6vY8+xUfv3KTGNUc91AWIxuTt5u8pJnvX0kLcvP7Qgjz9MteTqKXV3HH1dEPFyYphU5vdK
tcLTQO3jy+PyyVg7Z66/+9ADwpdJf8HR1ffiX3AQgwKfs5ljVPFeptQ4PDgOTidVyd7nrOJfibqd
7uYqjHOn35nRs4O4sBJBp4ReRMEet/phNJjxVe79FemuTiH1F3gJFEOOdaN/AZxOMOd+kMAv3C8I
al1fyEnEBHSPThWsu7mGIqh7y7XXKRaeWlt7QGnMz1EoxoTUIRE/FC0IZ/Xhd4Nb0SVKo81p9wO8
zK5artOJnLGY5emJhmXknc7QhD5RKIG1p/GfyKLreaOM/PLCcEFAKKAQDEiOb8aMx0vYm3razoT4
++N3vPVRgU+E6Xb9b+zJ1uttlycKm59ngtSmzLV+AYCE3xRylk1lvsZt+pqA6mq3DxKUlakcJH/Q
mu6LhY5/fp/WkbhW3pMiintN1PFQFITtgojOusMyxeYt6ISpXJ4OTTyqrK1KUfvmCynPuIu+9Dcz
fUwb0859R8G6XEFEP83mF3Dl8aeld1J5hC5MkXp1q7tdL4NuHLn5Xb7GWnpD582wvPGMahPlSIK5
6VrpY1n9vz8ZxtWgUHJ4wz5EKhUbe6v9TkFq89pFQu7gNP1Cxzl1dgdomOvEaN1zD/373H4I5A4c
boNh84fCZZRIVwOdUudYTTKWDap5wSaCPSJ/9VsgOeDlkif/u9yrrPqa65p0JRWSR/F3Qhygu4n6
5xiIVCIPkx3gHWo3UGmjZ1NXv9/CcyxXn4W/Ojdx8+VtMYMQcsJaji1oOiIa9z0Ba6VsBZZ3ecVs
9xYBbp/2D/kdqiTtNP/gQWwEI2wIabzpAi+fD+I1M0D5FFxFtKQxehkuNlucPeenRHRGY/+2mitY
TtaRkHgE6xwKmmagMplG/otpWRWhJLHwFjXosiFFKghvyVCKh2d1/n0ZjlLyK8XxUZ81YOEYDjO2
yataLAEgHpCcwrriMXC7LxXeT0g2wmfipuNQ2tppg7KWHi1k/aDkvKfWnSbnFYNDTO9C2LCQLMKC
1WaWPSoR68SXidNTDDMsAdoprtWoRvcENcgaUHr6/4zObWEqhM9KSc7Ycrr/zgMrhKHPhMDhsPFJ
hH7nyAyZ0DAn7W0ZYIIBqbrg6OkAxBPXTQI+QAxcENwd1H49z19Xl1fiQl5bJCaRUblhTAb2PHvF
r7Ozz8KbQIFbma0wGvIMMeJWQKl4a+VQZ3UaZRgm7FC1sBORt5N1M8tTIfTJ7V5qjLNgHZIH4Oa+
SEjc2Kb4cL+mCgerUK/RVFJGo3kTgve5FtvNF3zC3ySL4e1gduiJLEFkSlBUkhuCEbVyLkSmibFo
0EcMVFKkrjfx4QQ4EcR1Lsqx8aHcreKwHfBWdc78lb5ZYnw2cbpWBkNQELpMNPU9ZHel7Btrfld3
iHJ1IZPEAicwJTMLbcF+PLBUNRqstZdriWxfMGfXl/zviUBfXAn/Pl9xPeDjbsYMuexktl6p5yKo
K2pE0BnM1coxuLmpgP4xVBXERENcLcefMmGXvav8vLXPQfrHOiRMZ4xYUo1kUh9uCHweIz63ac1R
oNbqIyZEYlqVAjkbVa/rnmP0JmZM0W9rUiJb9SU2WnZ9Z3TjC5/jAYc6sELPD9oO92DQA4/vlEY9
CtL4SspemF6AQe150irvfHGdwq+A8DnfSKJw/JBHRx44OIq6t4ohsgmfD1+9UGCxXCXXwUM121iO
DhDVycajkWNCyalwRL7KN3onmPrjBUoc8MC2C7SvVj9G49LmvYc7tPrdfOXu/8vOAn8pOGuVqxbC
v8rHyDfB3IQEFOk/VENW+w8ZBa5H85v9a8J37fK24N0dRjofaDmtx/tEO294UN+U4qfpLzyop+hs
9TeisPeYn6htylOfRU3xYbW4LTgX7P0EKhBBMIWNo5Lz4kUp3jrvG8qWUkJu9/i6S1n+vm25Bvsb
iEQJqbBPIA+AK6YZaaSI/SwfSv6fnOinf1p0+inzKrWBYr0itkRauwsteW6sbD3RyB/NyhBNk8CY
o013NSLU8hTRjbkr9/GEFTH9+PNWhpX44UqZdZYB5u585zAM9yVZp861x1c4OvLrMdwJIcgt0c3g
eWdLB3rTLEWn3ms1rs2pzeRInf+huNxNX2HmnJzyejf3MARSZVa44Z4WQu7tT3XO3IfOY8JaK+e3
gouxWd8fB6N++TnRrr3F0B8MrbrUQrwQesvp62X0KBrfDJlcyZbHk02L+msbAOrsEBjvklawZ1wx
72BO9TK0E5IqBtdzVUOnwsBIasozr5vi4JVvPM/ZNlYfOFHvzOg0jN7N9OXGSvIvZw0Y0lkPpn9j
Bp2ETwu7VF/FY90bfc4Yp5GLg83Qlb5d/VeyJEbRrA6qEWVrtGE82viMhjEmLJZfxCfTXaZAz5p3
wDM9lwSaWrax8fQd7H4sn+0exntjwa6XlbjNQTy8aaV+zKiFo4TN88I9xQ87c5eEnKmqJ3qut36B
+TdRGjiVOAXxoVaI3EQNbNEUUtllXxIUOWbPQKJfRlUloibZ2I2qtPJl4eNlB71v2sPwkcTgBfRK
Yj9oP74mTtKIxmKiRBneUcsZJPkIBwRTYymDOSs8Nw08WjmZV5puzn1Gr7PgAFDWIbGD0nK2IXOL
/W+1w5lrTm4CLDDdY38XpILq8kPA0ZcJQxuYm8NjDZwPq0eu5virvMhuky4BBRqKLBCqa1WjF2UM
ki8l9wAFA4jz5WQ25tYRxZTJxFEcPPfFkY+smycuidyQzJwQy785J+mzyfps7Y7gMYBUnDWTqR+3
Ua2FfcfSCaUgWQYIadZ4K0cVRlfttwcMllP39VM8UxQsBABNJTGIrhJsTn+sjk/3SpgtVkoWsPtd
jDHcNQW0FPJtiEh6gjZmIK8TSO/YQNzpL786PfOngBvngdBUSbglULswz41t15uaVxdTX/Q7QzJZ
yKIc88QVGoTYBsPj6X4nc15P0jOkJTrdFObJIWGxd0AHhGM4ocrMK9t0FhfwxNCLY0ZHhmQH5OQx
MiaGMKcd99hSMX/wjrawEyAWoKkEIyXrIYmkpOuoUrH5LZ7WWyheCLHruxPLD+wWGKaOMOGbISyQ
JQP8gQV09yeoU7wsLYWyKF5L290xC2vh5KwmIRubKYunpUOPD1tEYRwbg0tUYVEJCced3JM69zXr
6WbfMJ69jNhiJpi1hqEfdOZY4WXMomA8RvG6LKRqWqsKkCKlxrvMSl/3iWt/R6KCynfwZz5kPj5Q
+Gzg3pXGRO13f6nau2775/DSMnPAh4KC/iyUDthIDhmZkCzwOQZg3W5sIwrn88b+QZMolV+t0dDS
8eI5Bp0p4rTAwevKrIhU9WSt2tnXB0VypicQzrp2X2WkH+9Xi8QfQbALSleWzNeyYd7DLSH0y/Qz
Biql2B0NyzI6VlOhRuTWMyD9cJ244YZlE8POyBIRITntRERRU8345v0MrrxFUUXsmzSSoBCAB1lC
cEV9wePIhn62042CaDrKa8mPobZcMq/KM9wg0OWGiLixVbYPCcWyysr1MJVHMUb/nTzEcaN228c1
0PV/Ocl7kESb35ZKDjHqFfb5GLt4pbwYxILcS4/reenRC8ZguokcXavPgmLjiKfzOw1pCVULTZOu
SBQmmb1eq8R/8FPfl4/aznKXuFJZ+5x1R/eJcFxNj0m4EFyxyOZ/QPrx7uJm+F6ImRnPKnwhWA67
o8/c5BDydfb87/7sVs4/CBYO8hkFE0LhiZe9p28TqRu39zMxw8BHJhYM6NJPu27Xu/OFMf2AsAYY
3U2R60vGKegADYqGsYayyB0q6/rJkX25ri9ZB+atJKwg6hxOjSS+7hO9PkSMrrl2rs995dGwP5f3
UW/g4qoG1LdQ1QtFBRTzYS3XZhAt5bgokVRBYjn4yfj9Gykl9u8TaVaUQ/+JR1K13Gek4HhMav1C
nhzyoC5V2sOBpBI/fakVp/QaRF7kmu6ZV9UbhH6HbjPxcv7dyaFY27WoVge2KR1EtT0oSyMCMUoK
Dzhot+CHz7OFuXtcFP/66WIHKxbrGnZ/IqcbuFMg17rChNSVo36TXsTmZCJGbi7mPeT/f5+NtwRV
uP54KxX8Rstq3aR4xPpW83bklBqCAznWIPyHCtC1P0d9SdZASqbVouUg2RNXuG2oFlcoR+/HGKl5
GOzjqZ2TXX0x5mqiEHBVH43hNpL001Hypv3iyftWleDjwbXVd85P0wZ+TDUQRzEf9zhvXL2JL2UA
2Gn702DG95ClbfgjguyHLP7vFqG+/9bLVsmk2DKHEYPDuZ9740mlKAoREFCNl1l4TCTeFuWIGdU+
/OOGDEnpF7E9QD1asRxFZADoziirsSz+O3hRefdY8rlodA8m4wnVP9t8plnYHJkmn+bjYyqyi+8L
AjaKbUvn6JxvgsneKaQMhymeCt1TbHk6jydsHnygzbRKcm4S6dJh9+qmM6ltz6+OEPzczVMbMJ+b
qMiLcAKrQROrB+5kn9xvrkBU+e4TVcQe3AE1OJwRsbjKAGr54/XD2hEPY9pUqHlEjv1FmBnZ36DI
HghxESfle7BShvCZ465uEKPDnd3fGiYFV/qWTFKGBlii4zVAH4+KXGm1tgzVwzNDiE6t0NUDourF
BcUt/MEGe1eZLVMYbfDguEK1oDudYSUZNWC72W3+VMO/z7wm/NsNbGF7LcdEzjjh2BSuVJX4u7C3
OQnsgKUuaGZRhUWQ4KyoJZUpns7trXDtkxl4e0H7zC4pEAKvBdbEEXRZO8y+iiiEcgfCj30Vcit4
wDARil/UO/9SZsA3nLR9IpoGthrZkMlaa0B+RRpLBqilN9KgXkkZcLuLJwfT8eBHoyLqffdFmtlp
mlNgKuPXCpet62/yIhg6c5A6ynCVXZ/2E1Cjxz1dbVnXiQK+HSmnrVuHrSOmJaAgIEdPnMDvAjvq
cr2Nxvg1+M1uUD62UGbl48qbZsXolqgBxhmT74mn6B20jbG7S2uS5cvuJurBnVQ/m6h6Z1X6kCHS
i6gJVv/8BZ08B7pNIn7om3nIYV4mVcEOozgtetgptrm3O0W1EhC6HZnZAtpuEjBZSCFE0v/BiEjM
L5keYXamMxNDfY5lsZ/V9PmZcX94CSu+CfWp4JFo/G1yf0xJFoa4tMEYJ5OgmJx5Y/rjmw2EmdEU
syCYg64OiZbt+YYtFOc9mVjbg2RP5dJB8WDLZIMcD2hSHtqLUV18JXf/xjQRZg+cF/k/6GK57yZd
TjZugGcCoheIeq9Ss24YMxo9p3LUSLUGvRZDCHXEj9osPml0kZcmBd9l9nX+oe0XP4eoeFoULOR5
GSzMJ3q/Ihql3ebFYs3jYUCjdDw1juPCdRfGLUx1gLRg9J+txaQolxbOCEToeL1W1muy4MyA4CFx
6bBYnRCRT5fz5FAVQ8Gw42aP+JcJsbxxHD2D7en8oOUHORvXZ/4mE2S2xzJb9KthGfbfanwEXxA8
FLCIaS1EN4U1OU9dNllbIExBrciGQKxrGGxbpmx4kgS8VaVHMGbd0bPk5/q6jGfkWJjiGA32v03X
JJ+k6IGUKl9mGYm38Dl1VSy6pqO9s2hLqwFAlf8S6Ae+3VSPi6WAgCcGO6X0WxGQa1NCnSUQJSGj
jWMm3dzx6HuXdw2ptC5CUFkjXm6sM8IxdZFSvaFd3K+IzK+Y7FGtvh+p7ixfDbyGP01i7yZFxF/g
co2tDmmb3JX7z8PXsQVwgD8pY1aWWst7ET4k2yPcLFkXXgpsC5rSfwSjC8DQcQCTgc6r+CVVV+S9
k55XNnQo5FmbW9sZ37Po60o8Yrw7nl0725vOJrJW22LKdE/yhYYI1hkz7JMfQ7Eeuaesf6fn+8Zv
Nn2ljJr5qxPl6PADBUVIxXP3fQy2iZ1GiDO2KIzrXh8kXaFKKGKJy3XnBPuvtQ8oo9n5zlTardHs
BSA5ZfyvCUbkvfIrEDN17lmmtnlvN8/FF3QR1JMAb4H4TtJUBdnTZ88gbzKw1u10jCmBVGi7Vj3G
JaVmKzGBEjwiZFZpwQdq88v0fgu8QSqyyjA2HTHuPb59E1RW/FAh7VLVOO0iIrBxBVo3lSjtWZTc
tshb8DIL3fL6XyYwxH+lmnYV0l5DB7O6z5ephyt2V90TmawjrhEQIhOYjnzzXWTJhv/0p0Xhefg6
lpSauKd/lWLwcz7sHpMXTGTjiwp5/w+Xc0NaN0zGGUn0OdaulxoGlornTBz/YnnZ/bXCMOEDtGAE
9UTUXyiUGjNuzQ6MEpsCwdRqqHqhrDzIlHdXxVQcMUQOCvZCHxOM1gUxCDy7gSzGZUcUMiet+8aW
RMgVXzyg4Yr9FMjdPjMX0o5FirY3J393V53+NjWmrG21M7/xuyoDH1Fh8+7umUoE87imm4l2TITO
MYKXeMf8i1WqPQQcR26jI1zTgLkNs6RSllV25XOyAHURkZ5F3JdLm2YJMFcFuXFvXIH3dwTclMCC
DcK8EuBwBiicoiqZJoN1BDKkmNd5PGP3X31aEBFYzii06DCcPI6fru374lX1AHHFPz32UvCRNcRl
9+UXWy6rEywlEu7gD6OYai7zkojLEC5IICsofXazQRzsKxd62IGtHjyfz92pHZHXfBDTTRH96VzC
5F0vCL8aNU/i577CNrhbSw4QlkNRxscdmyuPDv7Vdp01v/HrXasAUHemRY4/CbPKaqeqhsOtwTVR
GjCR2jvjceRU38R+krY3PrJCKJj04pAJbEcZED4B210ZeEBllpsTnjpoLN2d0bRtpAp3idtUd4dS
88R91KSDnCMUI1CsmAjz2gOIkTDrHJIORRcUy8cX+9nvWFLiunKTKMnJRPRmtpkx3iQfWLs1Priv
UvZCSthqbEToHMHzmPew21r6pytZLI92tJbUamHjj6U2XGUJgpwuV93Td8VfKtpQrUgtL7Ok92PG
MHCuha6eAC0OwmOMeMrGAXwFGW37Um+aC6h9GcDEr3d6z7fcLt3/2R8NUQpJpqtVehlLzQrEbFhw
BJGVzT1jmaKtTRp6PWULAkyoTtmtHkIwXtuwi1iKV0LUkWjjmtv2rXzHPPfBVO6ftqEo8o97sfm2
56hIHgfNW0Bx9LwODYA3H88mJFv7k6/If6VuuAcZWujW2nTXF1VzBPJlYPfl+g6Qk/qRbZaWs5Gw
pcTkw4VcWzY7OCaBYQDJhF80hoOvP8pCdm1jhzhrn/rtEsid81VcXNsNhHTs7Dm1RMmbDrfSmEU0
sTnZkCNph6WAGQcD6UTFtnLSzzMxbcR/nqxYpfQYKDcKvAuxiw3etTpiu+NYh4byUxE/hPeJXj/D
JkhaaNe4UukjfAHErVXqqMO1YtckC7gWXGCz/2ZybGsYBxE0WOAWzecjervd3IvWW23PkpGUvTa3
FdMDJD3Ut7A3bVSkHRjo6ugN2seYDkJIDRUn236uqvtok6d5cxjfKlaUHWghE0nbltKZlDg+CbbI
8be55kACU2ur1CbJexHZZZsYxEKNnbjG+jnE8A2HZniWlM2jpVjycO8xMay5yqSC1+FnZZ5P6JiF
undDQPeSjYHiyht74Dp/XKj0NNrpnc140Y4Wdy1DeAEWu6F7JGorhXgBaeILBd2mLQt47zA2pxV9
Vl+umrP/i8r24VxGwNsGsJuhxXXmmFKYmFZgF80g2nszxhe/DR+aQ1z2DaZf7IpciPEu1wf4I3QX
qsGaP4rctLSZtVAFpwnGFw8vvpylvw9/yK5jSVFjyB6dTmSvBP4M0nDaVMHaiZIsDTia6hDxVqf4
O2shHMEyAcShKuZ/gvn1bQMLT8KifYMNjGUjGnbBxX8iTgH2X2lcn0cMaT7LUon5YM7QS0ZL1oUN
dbQV801b4s6fl1waXCk8B6oAyGRiFX8Hg2pkaUFmK/1KW2wZSX6CFO+jRElacs5JNeSIpdz58nrm
OLQcYCRMVN3VkrG8d2GlJC7ARWW0PNWeW+gVotm415+wuip2jEGMakpgSRWL5aVBKatECBD1rubr
nsd2nfz4ahUb+ffpxy6GFS9EYZm3ETx3YT8BoF30AzoUJ3x14OOpwsAC6UWJVT9bq3SwOfJcAKGo
ffYbBZ8YCWgLjDsa4d5HBnyR2gz3eudtDkSxINgBKARdGnEUlava2d4HPbJUJ7H4FA7bLhYVN/Be
hK3skAh8NypTO2JUlcaoP22Zpgk7TBSTS05FpZ5838unY197Th8AqQOYuWUGKEEgMnygJ24dtqk/
wSzDv/aXUju1gLCoUlJ6Vq8cP7sJU4f/LHYIvNspZkYcAumGtTv3Bx1hr7I0uC7m0+i5gI7bBXtS
7e68x+x3HBrgmOFvLO95DAVuqv676Tcr+HsdxRauOY/Q9wnnwil8UX2+pIsWafA557T5YZ8Lbvd6
c58JO3qnrhX79H1zZI1Xm3oucSMsN8xuZR3phpHveIUJgfGFHL586ypBwzPX2AjRXINL11xFw/7Q
o+gImOV2h7qr/QftQqe61RFQw9uB7adWKLjg66nXFbcZoxLtxX+t+OTmPviI3LAwfIOltmjlphEp
Gcdh90INMC+we3P+kNy7cNKzOgVlBG3ZMT8EMykRukG3K+Q9xbenetj8ZF0oqcND1XT2pEHPyzp/
35k70MPkVhg8z7sAy6ERRZmCnchev0HDSmNY7ppxMn+4GQGQJRbc5raELDb/6YIJinUbtVjbxc89
mC2Tpj/3j1k0xWky3AAYL4rJJehWDIvty45svOjhCy/XKHhE1Ik9lQaICJ5FOb1o56jvCWIvj9dM
m3gE0ok8lKDDe/PLF8O2XB7v4krZDTbdaR4XtK5fYDmbMAMLU/qoHd+kz8w9NgqAosxLY3V5L15I
exVs/6nSFw74rKhBiPrZ5x1WlyEV+fjBggHbGhU06NAWETGbjHoJ/bd3MVTj8rdJs0N445BoqjXo
TQ/oW8yt7WHvgeYYuEQQNrvGqCS2s4XOUCptLnEl6sxyIxs72XX6FIebTA1FvGu6Do5J7ga4oHcD
xfMcPtXkqm2wz5FLqF1Z2Xied7y1UtcrQZA4ID+uhfNkl2DQ6BgOlBcBsPnF3aqmq7PqbIMXmnKX
7bdtdYLAdBf9L3gUXsKckTf2mjpQRPr8ZaLyhSJSdvOu6dal8XgVEU39uFoDsZP79BAbiR1JWf6n
/HUZ7H/ANhmuCzLNtn5t7cK8Z5pDe78b1wZ3fYR0hLGh03ilS3zDQOlUyhziIzITAM/G9LKXklSH
LJSZtfP3lbFd7/0e9VusysxZB0j8X1oqc7EkD3VM6Iu828vEDzXPYtVH8nT2dwjqliqGUNUGIPAg
abKD5FxNys+R8D8jiz/0EsdEgv1FvzSovXo+kURFdYqmw2kwdBwEt++8W6AyyXwT9EjFcbtV6RV9
55UMQreQDPliwvY72XGLNXsICnRKC6HzmMj24H05KObRLR+WeEEfDeB4h8QSNWRwilYuruGOdvNW
4tZCJcGHwyOZBxnFmmBHfkhQx6K80KLKMSYSkk+ywVczgmcou/PbpnBZnnElvOya02whU0A/+SJ3
r8NGi66PY93KlubuqkcqfxcK4UtjrAKkgi0aCrQg8uz0l10Ocq8Uysj9MMLwiDh/UKhNzi93jWFo
Ewbmae7qfXR1Z8WrAuWydawkyYVRJ8dzZl+RAtisSOBAr6vjfaazZgajosiDA7HpePavCZFUEqJR
hKL1Y6vBj4Q/dCuH4qEZst7pAoO7ye617FMsGC6UXodnGbA7Lby66EUKUyS5zVRCmbrAyC6tFdtS
aqlBeK6tJJEDFnlJcbq3rqKMqB/l/AP6T2elGHjmNXM1iqSMQpugF555wQ0Hn5sMKL4i8r+eGY8J
1IbiT9lRVbp7Gt6nATfbm82Dt2Kl1aFOl+apVLNEB1EhJujU5kaU+UkOcnJ0r2uBccNTPzSFN6dO
Hd+9LyySxBzPZvItEwh/ZkMNSp9kliZKhffMKmswoQLA0XAtee2SrWtwIpOiaR9cTwbnXoJWqU5J
lUXHStbIFBgSZKFm017TG/38hBKmxGtR7YUovvwKN/YxgQFZy3zxC8MYfg69ludAS4z//7KzCSMb
R6YT08QZJBWGRPqW8afjIRKNmBm2w97qUUhM90l/1NN1n6sMBFIrimCbeQVMiY/cZb//0AjIigSK
3XuyNre1Ny0YPNd15hR8JkLqajuE9zb6GzhHdXg+3GvXwTLuL4pQM6GUKKdqHxOWFSISBdYlIek4
Q2Nw7EDh2pg3jQjKNyURX8DCBecKD0TYnwKcLVzBuIs7ieekYhsFfRPOia3IjxsynykTcs/LxwHm
XpoGa5h8GNpMNeWGdmn/YtguooKzPmSSKSKDaSxh1j7uGe2nVK0h7mxJBVdlDRjvXHPS0hBLcBiv
Tdqsg3y+cZKKUh1ZVUagXe9LW75fH3peYCVbAsxRbuWZmbn3v7HAp9nd5Qj4M7/DS3qhsbMZBx/o
kxBBTPGBCkxOp75jnI5+mLmyWlBcq3t+QOQTQGoGqKkedL59sR8ls4Bt3+5I1OmlzOQEbvpftM8o
jsmPrMB36hOLPKtkNTYvKbdCJZocFLmCcafWrMRCVGoY+IPBenVhqcuWhfWUnfnH8wev0efdbcYE
RKQdY25I9oe/s8kFcn8sIl0O+sSnuVfDfm1B2aMlcvntEcZw118decXyZRzrr8arWt07oaG4DWsF
z5en/aIwmZ6RzmiAKK0jfAEzAW6R2+ZFsSi3IXT8HzAvHKWnaVug+WOZw+gi3zOek+AVEiSNm3Dd
YZ5LMnTrqV3rT827eUSbaQxbQaSLyCUrEzSIqu4cDvHfbyEkemKhGZGZrK/QSC/fMd6yt0nWCcyL
vyesrkDrF4LGWfgToexJs/VBfaStuQ3UvrfHuUHRHoGE2jZGrpLTjMSl8s6r+m7TXwe8vnZCkM5a
9vQdy56c4qHzxx8F1mwBayOjBc1jSJ5rijFxXR4QB6caAmc2U3sBpzDNxCNk3JwEZMQAyrqyXdDN
WWwzfhkf5jXommV9hdrMNnzA4gFob1odBAt398TSUFtFRsnVHOnsULUDz+GT0jl8R8dxwLPkSUMm
iPjtWo4kX6ONBxcn+3gcxze8lpPyFEbBUF7Okza45H7ezo8TGAvZzfg2UuESWKoneGntoCVt37Kz
+50k8aXq2PXgt42oiyhUIlDfTOhDTCaZQNHW6L6yoNKirGB0cA27UarWiXbIyP/yD0JocuQ6X+2H
Rl6oXzgSJHsEB5vaPmT7sNVr1JvjvfHkWvcx81a9RuAI8HnVsh6nkwZ1LA0cjUCvQRT2fKWphItQ
24e47Z+hknRo8jJGHA3a7883TfpXP057wcgyJxxV6YAQhNwHH2rcHSL2Faw7lNJVefkHkY2SwkwC
PAZII9mdnNmf5Q4JH5yVeovxiTJcKmQa57SueefDgi7Ea4fuH3bQecAW2tW0uqPoRaCzxNqeP4s3
h6ywrWNf+WCWt6c06ACFXrh5gs+iiXaY43rwOtDaVoOeRa66goeIk33/2sIgPnIUXQUZ4JMNH1Xh
R+bFWdRQBHV82k0bV2TsrBN45tJggfUXAZnJ+kGybVjWDQZAdWH3XD9mGIYp8EXjEWEq+GinTJ5Y
06YqXOd40BR6idasE8Vp5vK14hxM/KvipdHccXYfQ3R+pI62OnZLO5g4WKfQQbV5TaB53ku37ayT
jrL5LZVzQh0o4mPx6xL1EYGW+mlRX9gXN7bASxuzrHYcIFeOqVKQCjXnPMBxdh1wWySC3qr6M6z0
dryUUtUnu1BisD2v2m7VrCtwx4hUrgtq2mie2Exj17AmfG/Tbxarbtk35MN/tlxCw3+qFhIEWa5E
OL85PCPqhre9Y5yHt5WAVftikHjyJRAA/QPe1azpSwC7jBXP/DT9f3tFsaGLlvtIIWJ/1IHjjVR+
Iw2AI3rN0ha+TLWKJVDZ2y5W2Yxo8fyaRmNhqF+VBdcwpaB59IeHDbo4U9kQIZLOQUMDnqyWj7K9
6fzyQcR1y1y+acHJ3yPb+zRLSplQuksZmp/26U7h7SnI8QcQa8o0KgbHpvAPYvHC/tx16g3Pxy4K
HMbcy0Y3NF4ihcd5IJ9fVMZ2kPhh0esk2U2sDlVpDZbf7i0xrmsoxi0kMS7V+6ubl34xHEBR7Hdn
raSIyXyr9E9VA4Mj1rOqdGAy2g2brIOKJbEQa7FpDOwMmV7sKyH9LZWK0/JPl09fyOGgAUjhrU9N
a0brCAKsG/iBEdtmF3AeRdV2sB7bsT7gqYcdTnu3Z4S5wE+qJP12xKMjINH3TdOkLPIrAtenWoOi
JxzDKhD8ogVQZKnGNvrOaZ0VMyiysKXjH6gaUEz96yejn8O7/a8eWAZESP7/b61/BXidqJ3affDS
wnUyGNCiCdVI/lXWovSLiFj3VLp+x9azbykWRzxA/u7nEvmfEQjkYINyrPZCy8pK/kYRQ2f5H3ul
iUwWcGC3++mPWh8I5j1Z5uDDeTGDQDj7SGQc/CAIYJHDdEi3xnJj81AFGToRTyeyb7gtzH2vIF/Y
xKnK0ZX10A6jy+5MHPClKD8JpSIY8TQ+0GpapPRhe3F7Z5EdNQkzdnX7n4rQkNfg3WnrEz5uZDQE
bbgCnLbxahAELvYY5zD/RLAAaZxLvEuQcY65qHwMcVWpcLW4N+42MeFARaVgplcNCEJN0Ju1cHhU
vuhebn0RxNuxz58U1flUPMj6sCM2mQiaYqmrxIdrW/aIyOG4Dy3bAA505OnIAKuXg9rmY86+RPli
L8reiCqZ6YsKBjAQ92OegoxzxGLCe/YkIdMOw2+CGRHG0koVRwq1N/++wCnp7IPORnEI81s0yyQA
fVqka3DoO/44CYWPkWker1aZeG2IoTxxeQnmla1RVkA/8+QJ8kMKRu71W30AtPs2YEB2BmStWrhl
mdeOxU4h6h/R9P5RooPk2NDlK070m8bHCQyD0tSok7S9j2IxCV+zvPaf5DuJ3u5b8TCccVRRgj66
64rpW5rt5IduEEi8KTBqcOfWVZS0aZQ25p/nrovvdt7TPjXujyWCVDvSvw1TomEDtPq6e97icsnI
OUzAIwW+noOvXfn0NXpVXeH1G1shg16k3wrAvRAxW7+qxpvODtmvVHZs6xYkDaU8JGTy9SOq2W7A
otSaiuwGEbfFcwZVt84dU7yUTb98PNraxES4Xv0PVFXnu3JgeRd8XkKGUXmC5pi6Gbx4pb0dVQnv
Xw4X4Ajeh2sHkSmicXAW47iZRF5gCZNbLggqCwdFXImVHBhKj1SjOOI1Md1xEZDGgSuvXKKu/ANS
wIN6eNqXa2zGN/10fTQlm5s7gAuTJZxPzoAPFsZYCOjBH+/jvqMqou4BDqaiX5pNzRfLRYU1kwoq
uzBiBEN5N+GHzV1Z9xiSH4xuCi+Tq9qVCEZj87tZhjiFEkxNFAv0BfhV6Dhxg4Zna8f3g4joREXI
V7CVQW5BLCqJn7tW2qL8cpCKezlWyVSV86jiN0Y0twnbFdOhideaJaVMIQIqqL4JfWMrPwlLwvUP
wV6kELoHbVaZk5Uak6alufLvRON8AZILNzSsCX5g0uvJHa0tHJAUOpZvnoHwcQp0ygF+ES2DM5d4
EQPYavT8enBRsMfjQIJL9JMbY5n8G87OO2qkg90DXWGYDxfaBEGfH4BSQVpWmB/A8yp1l/oNuMh/
ue7iFlwmRzMlOOh3YVI8SxiG+395827YatKoSIFMh/EyjHpVGn9uQVn0NWhlKOPAV2GKDgIliTVg
Gny4tthnrYYmhlTzDdQIwDqoYJq6jUqN79PVk7esxOpwLNz7u27t82Kxh4Q01dgfUyrVJra6uMpT
hlkKw4Z11bONYL9n+eJll+UF0PADddJQcfg1s4p1eNepBL7NusXLU6Et0J72oS3Pa30yc3RheMvI
uOmh1KPpc9GjFkXH/FvGm7zb++uvNnnP/rJPNH2DApixejmIWV+ztrcC14mwFkHFwpmNgMb09hhc
8hTuGQm3xM2WPgJUIrkq4jXtfx9j4xgQZLLPV4K6coSFUumE0KIQwr8tYlBh23/bufsohzBJHCEk
RKeq1UgE9SmCtL5oWIGI1aNR0rjxbbidnDg5foZ8jmM8qXz+ZZoEngo2wxzdarNmDUg3I4+4rMo5
MhQkGrqzfYVX1BXdt22p3xF1LlUgNw9CgnFR6zultLvHsR3y6p8CrJsbXkIc7d4lFafZ8tePT86m
OW0F+eWxGSEY8mtaEedonGWPv2GOlcC7uJFSmdYc/IHuv4wdmYDalMuyJQLKh03IuQv9moEJmIv5
56RdaSolY377uSPl8vHIQuwyJCBYvg0PWCwzBhBQraW1z/YdclQGz3LpMUcNAtN5yeYyHYxoiEhU
qNOTfYImBHvvYLe2hQTGlVdp9kizLxS5A3vHhMq5ozOvRJNWYzvl37PjXIyHfy+X14sAQ5VmCy1b
R4WvaGoEgFDM//ZBD//yRwoWsoD6wZ9PCTlLuD/VfISM1VcDHxh4AtBJ3YBBuyN1GjUA/YhApQ2C
6QwLQjmuTJI4gp7m5V5Oe7Xupuw9sbi/WNA3iqBjseNgvle4bcdjle5HuBxjzqJxsrW2UxckYuGe
WZD7NntiZReEU8tAyd/mySqJ8oBlYzf5AC7t6joNiR4WgPfSFWG+dndKt7Q3fBY0mdBvcdqZ3yZV
/uROAYcE8E5ON5BcI8c71I5Z6TKrYjHhxnoRLHP/dz0b9DOQk64NlZVIy8TwJ4zgGd1NTKbCvP//
867qo/uCRN3c1a9SxEWfLuUyqz7E8T1gt0Gv0imca5Iq6O909QdJlgbQCiiss51Q72BNnBZNd2D2
xkfRnbXDmlCX/yCehx1hcN9NJrwbLWj6b/NU/EorBLZbrMauGe0LukYfuGiumbEDWwx5R+fW8kYZ
xt7Vt0jzETuPrHOscX8vtxTOxxaumWqRhXjLmMO4Yk2jaLnL7aAuZESanYKqBh8s5f7ZolcC9NcJ
nzBiY8JDVWFj4E8Jhgl/0PDYKiBz4GPNOPD/JFPM8LRC2+prCZMbFTCe7+1FD1WSSsSHu1yu1rnb
dOM1+6t2H9kamKsHzLZDfVAKOstUUUuY5Sm2z7KPgdsJq/Rl9FUm/3WDz7PRZE6smkpUYF30HErI
XwWiSPxds2KoEFg/2RUeUWUSw5x5SAW+8JkdqpD8eia511YN6CGP69sygPWSl7k/+wbrCYB7pzUa
s+pg4K/8M8wCk23x2q7b/W1uOBoSTMDqlCCPwa4LSaXhl8JU9R1OY+qXRmfM8zg/Jd9fC9jOTo/y
N8h5G633UA4qO1e5izL+1VUHj6O6Pw9MDY9MuLXPICRP+PTfAtrUq6Xbo85v2zpt50yxYpipFK8s
pB/4u/z7b05ruAeIxyKTRANITUG9LwPfKr4fJ/jY1vO8vkwEZdMaMueAO8Gxm0i01pnzpK4hiEWg
VkauAKerKjKIpRsqXyJVgx5Y1bJPGDwj3l+rk1XJ38oARMA+yCWGfwdVW7A12nuHMrtj84ixu1Zz
d4wszyyL37j4W2uj2XsJUFk5FuVysWXw5phbBXXhjlAm8n9FB26ab/NDJUs540/b06HR8+XUQzP+
aqdb9zPz1N5xTIFkTAaAcUTR7+YeT451uBvfCTChOh9fXhshL4oLLi8ufbVeNeXlCHRRDaQ1TZyw
0HWUpmgrEJOJy531Lr18gbB/VC8hQ1239f0pHM77sJo8Ysqjw+aI39tVfjNJlQ6Ys8UuB+SfaNaG
TTnuUR7l+tjhsy/tGQmIqd8N8ny88tzkOyWUKJtN/RJCXPZfHQopVmgq+jnIm4NZp0B00hDyJiRj
tL61hbuBNW9qjOCJtsgf27xuLgcqIOHBw+u8iq6RSy04J2AJLX9e4DP2FZn62EFyUC1kCXEF3vP5
kQDUVKOw55V1Ex49H0RPwqidoB0xybfmFagewbNYnJ+ZRQh//gtCguesiB7TfPFwQ0NrOjQceC6b
M6upa7AHi3Acuof5ag7u+F1gr/wNulDI9atyqn4R+gF2OrmxesPWhhzHfKOUyqWooW6yRShjKEiP
cli385/Q0xdsrNAsvBq6/v3rNn4l5v8qKC8xrAuGZFb07NZqubgnYl0eUfK5P0OFVpARKac64lbG
5Tk57Obvm/wpvQBALayisT5PvpGSOxSH6qFbNi929w9DZCBe0CunCmsIQIM79fD3hhcOdvR7POKI
Jlzw02rvu4sibcA8mKHfmMU347HsxdjPmWTzjw4jqmkWHb/x9ps/nf0WfJCZ0YEYcG86u+0i31ng
iDoAjXQO21bWal2EFlfOObP1ANKU+iy0VdonCMeU+LS2vCD00PzqVP0VEQdYUtUHQGFuMINFwme5
jceiGDe/QIl+RRdif187MMOXBUiBPasvFVnYNOQ0tRd/VI1BmGKamTnoj1wIPjEuksd9MYYFLYXL
bPVMrqS2zauwf5eTHcExHLm6baHQy22cEjcwyPL1GQli6JYl3BuIjd+SfifruMQ3m8G6OVFcC7Sj
iId5uaRKRLG5fTzXIxMaBteKgIDwpLKQYq59PQc14rpehPeZraH1E5M7ABBB0dAvpEKbPhYIHsza
puLKjI34Glw7dXpYnrQu4TtFyhF8/lVyQQnFx/2rDR5QFtJpoCWP324+CTjuOZgHhRFSO+Oqjjvs
0biyan0Ci8uBciLNrKQ8ZppDxTUjXaKexbrtqYccUaUqncwulAhnQkMWCEIBwuv4zmPEBSvgPuAs
DS8BosnvP13ZbVb/PvfM3wOiRedLK4b/faK8+ou+ph8nyP4aanUD5xQRTHQ/j296ULWUNn9VItd8
9d3bpQgxYzp0DsLMQklyywoRN1mSy3nIE2uieir34/8MK8eIrRM3sqPRa0FfM+cFv8ECs0yi51rH
FArab9MonxgYIyq78g8pC8FnlLUEoTx8zNRdy1t2CPvW9RYaudBB4N8B6grx1T/IlbPNNEFXDmK5
DgjTqdJuQcqZ1D7KfFDFgHUNWj7pnnF53rwVvp/wzBmWzCfMEEGHL3H/ZMm+K443XB353LE/X2lB
G+TVVBC5H8rdGg5MkQF5fWmFIgIHANuAQP1eGsfJgJx8I0BXFVV05PnngKOcCCXKNZErqLxPmS+P
AwrpAcJ876ftnlSQaZdxZkOO9zQvtlMrBbOAxUceHOuEGv1K+WisTAtveA2f869hy4fS6nGSgLV9
pveCCyN+huG9eYIkCIbujG9yaCxf5DOwqXXRe+UDxqPqYleoQ9HMvNxUReIRCKlYBGv38UjTbYTb
lgYHt2RdHnnRpNwep0VXK9YVr9n8RCkrYpxE8WpWgKJsU5exJRVZ+TqxRzVP4gMRJUhW3GBSj82d
k3y3AY2vvtUMrcaiSdc2r/KciQbytT5Ur7BY4Z+6haVfKfDzn+wq9X6lxf81h8BWvLF0Gg6vxvZi
NcSrRxDFQ6Xq4u7pXordNjkq3/seZPVE8m0pKacnjMdjykw37/XGASYdMMS8A0MHGhXU/e1dCvJF
bELpkeuoHUVRGoB7txWATAKJW0xSjSt3uiQQ+P4ERXAzeAv3KFg5Egk3ieDlcaxuNlcyyOmYI9Jj
e91ozMBrhM/3iydLNBpCCPWq4YQZp+n15QOAsbxWDzj/GbuIncLBeHBsTDZtuLAMh688/w/h2O33
Um6cjye3tMZGpZetoNzDYFHZvnrEsICGCwuufSIxBS6LwM4/Olc67lfybOE/qAm/ptbx+8gsKJzV
hsjXfXIG8hKNifZRzQOWMQqnheV/wppWlFmgMU+J4Ny4lJBLW2cGWznrGJfoKXn1PnSCTfhJCrhF
Ee+dzZSHhRUjUG6cFVkMDi/mwgjbE54G55CIILlm9ocVPce6eCyiEYTEMtqn0XuqmhqXDlK8FybE
pV2MGUuaYce0VjYHlnnePTbQTcQ14Sbyi81hKKtmtDMXhRBt3dbhYL6PrwiWdWSeldl3w/ePYG0m
Mt21wnYPcD0AX/wmdSJ7JjlHaJICtZ8I17itzm/+lFfegNy+id2huPNh4718FRdkcmzCvzgeSec/
dusbiP83iJsSmsB9GeNNHYRzOCivt/oSQapWm4UnUl5GE70h4DIo7Jg7JRc0mZxTPrNwf797Rehl
ULDDaijmm/9kMbkpNTiYT4f5kfsFjR/AEU3/FvxjyqtW+7s25SQwsmk5OhegosuDH3kWyLIDf+Nb
yjK9OkdNqRNhImfJoJP2Bm+KQCNQm7+OVFnMWIjMpXUQYTEx8Dm9hOmsn4Pl84vTMEN6Tndsv12Q
TPmW86eXsiAuFhPwGfMAwE/QzgxNHrnIdGJVIGyH8cKL1hkUJrSzJWBldJL94nRWtafU4BRPQlwX
yAEtPjs1LLVf9rdlEToeD0fmv1XdTez7KbeiV9H6s4w/wE7PcqvGnVFzW3CuYN//lZmnlUElgAYr
23XtVY27sXFyqUX7a5ImgQVi30kNJfbSqnFEPn62IY6yYcvA5VYoOiRNuvQcHx1VPl3V2f7IzSxo
/VDzJpSk/dKfulOoKqPxQ4R6nK3VNVp++nJmgondk9AkIw9RNGMJMpNSH9HlG2IqYLYxpgbx8vQ3
H/kJ7TO2a+Q8q1gqr8QLs1wWMc6nXh/Qm1g4IyERxT/WWn+MtgWslKUnoPJ9Zqy3ZYNrzqLuiQam
/lhs2v6UdpFkRzSMg3plkgfXofBdy8pp3xeSMhP8VvheZsjBI2lY/Jz4C72b/qYhN3Yc1M3dckJP
MT5zqh6dTwS27GerEEUGK+JPM+F1EVzHygMxjYSxNE4MGnNio82iAMaOSugC5r9RX9/fWEJ5soj3
keDdUOUSXx0vwbT3pA3ow98uJ3vTZN4SnAuGGUbHiQqzU7td0NKoKDwTRzdBCckjkf0Iz4GihjNR
SZKZjDEQ+S7XMUjtOPDYaFiIU1O/J1Tw/nDB2axLTRyQhwDLsjQcXrttM2l6L+FrFVlAMRy6zyNs
qfOpeyHB0yryzdRqWeEedksTZDVdOtCTgicAmY0LNY2s4UizsNqPwu53SZdJLJ6hqD0bfdXxef7h
ys/fALVLdJPG1k158yg3f5vfXXx7CkE5b/pUf3ugdLI0zTm/o7G4AxRtFD2+Z1kZnnxopkHOVqIj
PokeDbEaaXtJULsIa90eiR/2camoga9jay1FU5rH1oo5GmsSJOFiSXlcIrmbyXA6eOtBfYLvlQlR
z002Nm6Q9Y7vcsLYUxIKjDx4vhseRxoWoGN8CWVoih/6R3JK1/6kNsnPPodJWovmJ+l847Do6BpG
/kqVewnhZjR7YTnsQ6aBB07ymm+pVadhTismFpzXsXcFlq8oL+5qV4F8o2WB1a8llkXSVNhikTc+
M40VKaWEvhqyyWaDP7lMemCGTmSG9b1xTatj7ebALfbYtTAa3Z7SLh1olIDl7ReRtRf8e3QoWfKU
re121uoZ/PupuqjnoCzFskrA9amTiRjgIYnuGk2o4OrNY4b0FFL5jI4wYYYMtlvutweSLE4y/q/X
QeBfGJQ0fp/hB/7Hy+FzX1t7ixZQTIOBur9hNSM2msJA6YH1QM4mxVdp0O50vfaObN2a51pjQ8qr
yR9CD3xwO6XYUCU4Rrrm5S/rEm/Lemo/qdeq6e9TiREe704NiekUEDVqGcGtNURegGFVu1R2z6XH
50gEtjjJE0wCfPYnoW7fyl8qem76YkniS/OGh0XlVwwkq1Ixwr0pn21LVOjb8xWy2gbEeF7sQ8us
GDB+qVoK99ZHSN4Jmo+2MHhAw9Q5ZC0gli6VPAjtoKPTeHmc1z6SQ22hvq65jLghpvlXRujbjLAB
cCJ/cuC4M56Kk7a5agEoG9m2cpwGDiN0fLJHzguCjQnhvYQC7cyPxntRJfBxAHnNjNHi9vX83pD5
aPHGq9Drl4ginAn/VE9KD2Vyj9y0ejO0pSUav0dGI6oxFq7niHFriQjDKmAR6B3npW04HwjLLZbT
yVww2b6GhPnq928DQAJlhh8wj85F+N4WWuh+KdyYmUubczis4oSpm96vi4brWh8za3o12HXCB7JD
1JoJ69K/mZtQYUAsLkH47yLxkuzVHwyC+CLInyxnS4ggoTIDodFmdw7ElhTAOpXhJWVJCHxeAjn/
pCE0dkSdF/Wv3Ku9etZlYMR+7NqZccNQV53oUS87semfSbdDupdLByabmDxbFLc9D5iPGyiI45DY
zoNRILJ3yT4G8K+qu+/FocR68POX4RyUgK8v5toDF+xCRLcSH05rptcVHLjC0OtBJkl3XgUdbsvu
q72Q+5Yi2YJYiTqdqb9DXBuerWY4VP6tb/qccRH+IAvGJOTRo1niYnIMYWCQ2/tc9tUZsX3fiivH
4DpcDSOzLhMg4xKVWffv7ypHjll2B3ZqzWEHPCPQ4lCFHAt20CN7eXj00UF9FfCJ1CK/OYcLOI/J
XaXPORBZQZl+AV5lfyKyx2GNKswgrp3aoMZyT18IwbLkiLynaoDNNwsARy/RqiM9bNlcLpQjbgvt
Isgo5ImIg3w6Fu4lzs0or1W6YT6ou+1N+2HwvBUqf+0XXZ7hG8B16eglW4ept6TTrEQuAtH1tFhq
F6PIIhmPkPmZiB1kXGdoJge639D7svR4kLw3hassdBryy7OW5u9dvrTSsnjstXJMuEIEmKbko0OY
EdXiQnZuaguSc/kBsfY823F+pq4fqRVe71sYlQwJQ5BQhRa4hbSw6HBV9WKFwAcwKKmF4kzgBBoc
1U5NTPgY0MS9E3MzhHVIWfphFqW2LTEw9h+QT0TsAaDcCCHd+a3IeUmOXEUALidKR43wxvHLsOu6
ZoS4r7w3B4ms4ftZqNOCeJg8tT2S+dgnJmJ37gLiNiVhu5oVrdNVFbH5xhmHeQfVN7t2fgjZizOx
J/ySAbA98r5kg/9ounX8PhTMe9JxIjINb75Xc0sDupj486oaQJu8rgKtusE0E8r7qB/TI/qi2ARz
j4i1Tkk4w6xzilwzoA1Va/vDpQ81hKTjODp9cKwu0G8wiVdMXpHD65W5v9ey9jvgawKvpyXtwjWL
nZgWQNt2eExCSlbttcbL9LYfJqTE3pxiexYno2Cszp/J6L6Q7Nr/ML9nf9wFTwA6CAqwTvcNhXi9
hgkgAVgKTk7Zm2XG5zZoqmD6tsgAshdReQBC4+FL6b0luURUI7rpCsB7ZBE1IBwtdleWmToIZbYq
0kXFp99bFHNIqKO00guOamLNs8C7RWvKnJ4ESzHXiKwuzqMg1bhlcUqkE35oHvfakDVIKGji/0qn
pGGYLbJnl5rh3WTIkXfrXnAIVx9emgPuSnjV4a//f2hSzVMI78ApfSjZ/QxtxU9oFzhXmVfxNvXb
jcsOMfgHD6JxeQp94hBsiOctNNtLKLCFBGzCTw+NqMdNNqEboqbD65K86i2Gu0PWeu+e7z/sCCfs
STC2vLJHAHYsILY5vhuZs+qZ3+akyyuXytvF562YeFwOugL0g1VosID/MeSBY6qILYGAL8KZrktj
3pp1ZHW3Qq1Kd6FgaomXXlVYFa0UOVC9Ek6Dz079WcTUlPSoIdIctGkLLAZD64gsyVsL1Y1FQRYe
htecKAEaGsDySn9SBIRecAFMag46yRUh6c8fW2+Z/sU/aLhW0dXtqmfXagPhvgqW2wK/YKtTAm6R
fuSPuItDUB+6PRCZE3l8w+ly6RalBQyH6ROTZvRfkE+n9i3V4dmzccJupxzeqKphtVE+IFOyvLS4
feXutV/2I8X0VhBfR66sU8Y6UmrFviRu1KkBrYrT6Rv2jfbFyErpHL+NYsVr+PbmvYgtCGCnq6Py
yp/9+CnPSUsLTFmUf96Wfnb8+m0pMlVeHS+PJq2Q/GNF4cnPSBL6E7K5r2clOqt9SZXQ6oWdoxP8
4/8drYIzbQdLufkupvLZIhGeFSZ9KNQ1QitkMYQeoGxAEXyyssRvcV/AAGlumUvnbVS56UdRHn26
D+Ed/RMHyG3UUhXHCdzyixxRbjiEAfIsA0Ian+TSVd2Ug9bD9D8QMXzhDsys8SdkkNaY9N4FboDO
qOMXxa+WKpgPR1yyEcNVN+wETSKFbxLt1N39Otwxl8V2HSgA1Ow+edOB9fdgOSz1bJJL7aOgX/Q/
Wq042XJcwz9jbz89DCUFLkQJ7aaz2O90NoEjC/IMOO9ehHSa52U6DnEDo+AxMWhVToBNNZjsHWhi
PdLoO7EAlcJKb5VnNCTW1BbvZRsEqHrnFZdD24l/T644HJa47U88WO6jR8UrKZ/JVN1np995hSzE
y1guZEFv2YB836/2Cdv8w931DCk/OP9cMhx66hY2QBIOs2PI+KKsfNuso2/Zw/E3lLGaKzDWH9nG
16yqUqgJT/WvAGHjHRLJmXOWBfLNIvTIIdMOJ+8L36gatEzv7t5Qs9vVqiJ97w1tCxld5nP+7Lrx
a4m63swCKHgy3F4F1CHw8KHIm+ZFTE9dLhWRScooHYXX/ylHHUWqSfCeNNF9vqSX9y+TXD54shkX
mHeRRFFAoJkTj/O0lryPULh83L9HnVlDt29pw5Sa8Q0lWfYmmQu8kH+ljeVtWvbpJfrYJwvJ1oTW
ZWm7qDj7WJ82raxzMiGOsc/vVPP/7uhGJx556Grb4r5Vu3+gyhzYyranKzgJVf6Ts6Yb6WQ2IE51
lZZvfET5fSC/HFv3OX5byB6385mYjzGlGeYr/FYxK4eU+PAfOPQvD+5bUBaqyPLqjNeD8z6Amfxg
y11b46AgX16yTeLQfj+JN2X3L0vzLPtF1/47j5pa1L3bEDnuKMc7NqnkwNhnmg0sAcbY0rgG1xfy
MQaW2ziyzwWCzgo0I7fwc6gYUviCM9HScLZ3YZS+z3cFiws00poCXc48iX4Qiqo4DKt+ChyTipAg
WFocjLKzr9eE4s7BA09WLIpLEmQu/t8PW6GUeHAmfExjemgd+fXcHoKmzcO5RHcsjTuOEInGhcy9
zrnxdyHfw6g/hHbtbB++Wb5vHkily6Oav2I8beZsCmufzt+LSJHjUbpc8diT26nnQ8ZxgXvQzmE+
8dxEzIzbYZkl/fFquMizqVlZMU7UpIefBjDqgM/ua0D4GByH7CHkePSS6VAbQaERi42m7TQeOBNo
ZnmBmIpSDKcyDixbv3yUBSCexbsNa1dwMt3QxDFtumB+xyNTWAos2+/QOK84DPW/kAxaCvAiGKj7
6V5ZSuTYUtWBIeB9FyMJV99H+p9psvV+3/iWSQs9DbsPEPoiod/R6mDM1Qu7z9SaYq0M5K+vbqxD
BIjvHs/ByswBTSosnUfHbsnSeD9IdAMVTTJOroJxE+/ylv+UP7LoCIMOMWeJO30xGC5nPVNAG6TT
6oH1FSEsLjhMvNDKqyFHis8DOEir7zhzUu7kFPZuonkSRvQR1NhwkyXFORrEx5Lhv0/cr6aKClkQ
TQmL8Gr+2DUcgnNpjYSOaOhGCtiACYG7Pg6k6smbXqT+Aa08/bUqopE8KSB24kVM/KqCMfcJ5+Kx
Y/0JJ7C9q+xTDisL8Q+MlB6bAQ94wgsEfesoZ1qsRQrRWF4OR5nAR5JnrOTZNYt96cEoqexT0/Gc
TAqdt3hvJakQ3vU9UK/PDJu+5JLEydY7g3eIvfKx45JpBSAaY8R1xXvmiKR4oY02ymTQRgl7UXst
abrmuwp8ZdoQBQA7POggb57LVf9wHvgQjESSSB6p2WDHEmUSbV4c8mSDdMefBUlil6xowYHBSB8g
muosH3uNkNhV/M8eCtC3dNOqvrmgG4XQqfz3Ocn6ZhMNZVz/jvvHTrBdcwVZT/7CiH2wDgD1bG1M
8ErY1OsC86IavwH+S1Fs1VCjNBBGpN/5x6MONt6m9jDhNbZpR66HMTnjYnN82RhUMFUQ7wRUzqvX
k/9VVVr01n97oGc834vYxfq+jUJHgaqGRWRGo+vPr87ldM6QqlbwJFZ4aDKbYhYLFV4eex/KfSca
fn/z+NSwT4/CZaYs+aK1WiH4RSDlzPPK/c81DvSX/LaTWuFLbl3twn5MvwKfI3mVfphUBdGS+bL8
1J58qRZQ3rAHTKfjQreDgJ6oDjVGJdzPJWroeSGEKlZaLpE9YZgc7gVW18pPHYSWGyQVneTxXLU0
RQz0YWztkOdEHEzMcoj9uCkQkfasWqeKLf6Rvycc7nBe7/C25EnymH5heOCAokyJRx9/W+L80Nmx
q20i0nD71azw4T+rEGuOm+4zD+KT6HU7B1kvo5O7zg4LiwJlett1qwm8jkUz+VHdbe4KaGQdpR/2
FQRi7Pm5L2I0j/Xpc6GorkSZhegG/HSVglQlCMK+UhUS/pSnxrCgJeIA1V1cESt8AnpciC6zEgAI
FFA5Y/CYj4+kM3MZocZ/esPerwEwd8eRestC4GSOIl+SrOIlhUFmQwWj018NkmACsbrCAVUCmkMK
xX7sEBzCHqEuOVmtZvnxuE3hBD2gzYWZBdjn2691H3ZYeP/gAWvrT3gyqVsFevCKEWcGConGvmYY
ELzOJiG0wm/xttBusIxGEuCp2+TMud8l5/ay/ulx0gXQetDPDnTVJ6hfdIh+NNPl63M8OhIqmzmM
PYtnZyvjPMRyEN+Nb3uSmKuiP/gV4NdvqR5/I+nEv/e55yxmi8boeQSpurX7zi52bn+rA3cHXGfJ
WbjFWWIt9vNDz5Q6Kt2ffaEEHpswJs6j08WInIH9FGDXcOVg57/cdU6tfZZeoePAH71i4Esegim2
hN8xJ5iqYv/trvtViYdZn/S8N5AOPw93v0maf0ZB7aZmVN4kTndTZoyj1xdB92E+q6w2Tz2VLHov
Ie+lDG0QW8zDxaF60tDna496vSM6Vlzr1lRKQ+leyR60AuLcHDgE1UcH4/SHAd/SYduMq3YN2O5t
xko4z4t0eHdhn7sQubM32xzz1jd06ZTFVEkeiSfwHy7wEKDsyXAbv19Ore2eZbwLAo0itUhO+dn9
uTqijiY/t4lP1Qd0+AOHfXFL+udqqYa5GeZ4TlIYEkW4JoEMCjIRDply6Ctf9ichFh6/3k8tBG2D
LC+Px4Z0aJ8/dK+9wq7u5hVBH9vqMTf6BMxQlcA1U1Z3gb6ClEHptVZiNwmTkl1UzL7LxWVHgByg
SKyopE0ZiAg38xtUJEdng5zJhC5VB3BY6n3VY5821/qtUExk8tw+n8lbRqkWZcBQxuAQCMRiNnZA
j3ddWwjqGApZ6YVVXPsopYk4xt8CEjJbxJdObPLZpE4yBRHdw2KWxQT2cbnew/ZUWju5ykjPUKio
dicMKPjTquNkNsMv0dG1XVX8+9D8vodsYSwMzn06Sx4olgGE5rqwtHEW3x0b+knjTUHfHzVPG/jj
DaPXFgy2PE28o7sJFfEktJHVDn1caT915gXr98qmextJPUr7puJiGzZG/4mpQ0YfKSpCZ+sj/oWN
Ie8URmgJVXHuCEpQcexTLtyfid5DiuSmOdFOgq4m5Z1DBFV5AQq3r7sMNSiOGg6YIY7KqdPfNQS1
Ij/yeFJpoCIa0Ilsc2AQ266b8f71767pRyF1fblyOJUjx2SgGGug6YwH06X1z8ujdGCCvY7tw9Ra
nsdZxBimGmlTFD8Oe1alETFL9kf0f8H6OR9vTKpF5cZmm1Rgt6LDptx0Y42YBAbGmJ5FIy4Gmb3Y
k+sjniuqfDsRlqKiiFUGz8l+SlZgHh79YDopz6g1dLNrHJ1uk3CvnHOTi+glU8T0LcocVVZmgXPA
26U2IOy9X7TkQ7C7MCiXsUBGd5za35fuKc5KzNatsnGASJyEpYYmR1SylwHzXPzDmP6Erm4/zfEG
nQpwuw75pLwWkm56paZaajD1gjIfxLFBVphfy0lBci61ufhH/wt/zrQQzAgqsR+2GVtemFVe/fu7
sXyh4MTzdVsEwdN20u+lYFjWo2X1mfQKenSilW8LY6WPfnjuCatAplvBoBFXSD1o647wl+Wh4TSy
gX5yInQBSOYeYXNdNcXBTmF5xqh0uM7CqKtYcMv2TJXwkP1GesCVMDgg/YqNaDj1VB9v6JMalkan
9DvRItN2Uiofj8d5vxrQqmTWRJaxTGBSlyJIbrgPERAwfOwIrTXqAooacwlLxKv677GvwfGFE/UW
Yljph7ERLnJ7DOuDH/zApJJLJWwNkCbOAgGLvU3DauO4O9qIOpmSjK1y7YsV5jmcEiIm7yXBR1gr
iv+9olg++SkF8yHj3dQkgTSMDZanp3FkrVF2Ox2QbXWhWQdbfK40z8OvZ6mP6MbFvoFEY8Ry7W1M
bfs/VlUs6+ZM5NQpdPgKD5q4E/QEvoSQZlBREmh8tX9qV1273wd2QBERLxFQq9QV0DDHg4TCy2Y3
XTDPOaxc0xbJm6/mqoy6/CGaqJSagjW/zi64N/koFTVrA1oZclOEaWHV8LLaZEhSGL7HcFS0K9bD
ONHwfVsKrHH9tX0xAInAdxSSkVgXbDVpyolVe0pVBjPo9ziRATIJ2iAOB1J/f1dLg8dr5qZrkeFi
lMEffdVluaQEcQACXrsz+/fJFCWLbsfTdtdBJ2uByhyJKpamYeb4zRQ2c8QaEZ6/5qXE5sjk2J2p
nJs6twlkaDAeTTfKcFGF37UpWtEl+EkaUrwQejb4OJRqhpVwwuJhx8ZdwEiy0MLCXdrnQ1PoAnz3
U3X5KBJDjw06aTSAXKKGOALdkkq9vbirJUqw9qw8WpBAsMvsi8lcO543Au3FtWrBVsjje/EQUw8M
RFLXV13G/3WklbPAS73UAj+InjVR1b0lPCGJJvSYZx6ky/XBEw+PlE2reMnwoDq8H6nwXoVkdIBr
CzXcBHLuUXUhHs50QvJdprAWOYR17BxAhvXdv9qwaIKO0e03rkeNH45Ws9LhPMKdX+omJ6kmr82y
JklEmyux0bAj0WLKnxX9WocRUhmrDoBmoiFzOR5WGfyrij5cpBwAOW+nW51Y8WM/nsSCX2hk9ybU
6lIF2n4FA5C8rTW7CLA5/jflwS0nRL6mXCl+jEml3dft9HmcmseAQ8v+5B6Em2vr8DXNW5rV6JSc
QfVy/UMkEWliBiZ75uIPAKVQSmc0byIm0jZzUnvUX/aVxtD+EeXn+I18Wld6nv7boQplPWjZh4iZ
u63HItdxXhZHcbTt2CcCZGLLEdkBnRTOiszpbGHfOErTVqk6gXu9kW7QPZKZOS0s/vSsF+S4lo+X
Tv0N86V2m3NLZGNbz9Al8QqJbKLmhnUIjVfWYGseNoqi654tRFJQE+clf8Y9+8u5kt9skSGb01Cf
QkbIw5jt98qCi2JY0wVxz0MMRZIgGBrtbsUrPulTTQcHw+25nieCFt6F7CkRrf1H+reGDOOQlhfP
KIA3W06yT4JOl8tJZdg/Pw4/CJHf23Y/elaBmpTSEjRIa4ElxErZctjgR8ElfO7j2QU/U6jqj5Ch
Kht7+TceDVEz6dOZJaTzMclD4D+EeJIizTLgJOZU1Wj7S3DDHE3w0bEcaZVkzOCBZHCoPV9qlXKO
20HWbCfyepiu/+boMksa51DDuU8RTnidu84itQR8h4ugNtshOYZc3qfo8rvgDV2P0SpOdXeDkTUg
QTZxZ8XJjl1MT4dNfkNNq4RoViA9VcFbQu97dpmKMdwZyDOxW4BEKQCKJtlucJ5SSpbfCVYCjGhl
PJrtvnvNfl9UfLsM7cCGPrFoIUE3ta97QdP+piSafi2q+F4jXo/nhkes9QyHSR1tsRVDsXLsFKLN
P1D1QJG/95EzKh+Yc+ShgxE6aJudbNZg8//nKVa4/MfsQmj2tcAImL2qiU0PAS9tfcKlkpW4sT7O
o/2yFogiyAP+af0jLbFGjbrFkMZqn8phKM2SRezDOXV3KrXRfQZO0C6X7EmBVOVZUlLaVR2vtd7d
45iz20eH4wyzkwKyNGPkFwY2HWEm0h/SZEbTTpMQzKqVJzA6/1R3O0utV/QN5bB+hJIdOdvyZgfj
a/BHdfY9kNGKxQuzBc97TjMdDZUQ3hDqhf3aLQEjHcOwJPwPz9Zdi/IvFXCwgTgjt5rlxNWhfg2U
fX1TvwB5QBuofrhWg6VHGY/REKjTv247OIl1iT5WuRTdcFzBGfIoAU+1zN3IrVZtQ4Z9xxzzLyuR
hvhbq7rEJdp+Q8UlDENP28iVxCfxl/syS3hx3EshPO2s6iDYLrzPQbcbH2W2fserksQWEACLBEPd
bFPsLJFWdunXsOdJ+6upCnLjL7+EmrcNJdi8piLMc0E6vnhoiwLA1HO7Ba5voF6zSXDh9dpk1syn
PiqPo/KAG0y1SayvPgrHqDaL25tUI0wHk14u907yfkV23dhH35MRkmzXs9Iji4/1+hQ1+6+da0iW
SL6flvvtk/2ZUS7XDJN+2HUXUTOiNaXK2/BCLREhXyiqoOISaUGvY8X83N59cRNAmDxfAFGW1TZj
nBDsQkODedRc3hxwC25jUb2SRZ8oT82H9SzdOQBpGkkREaXIqTLKh0j/WM/8h/kck9YzXUTFzVg4
CoZBwDyTpS7r4rg6Z5an3QU5uLJ1N+RlNyFmTz74rGklb5Uf1JM9+RLfgbJt1/72yfdXoz3LvxZU
oSP/LVmUkzPU9178xzS1kxYI6Khn0rakqm/xaqgl2W4uGkFhZL/arVhAxfPWiboirXLEvi6SjHEp
xGl8IPZAgJgaY0qNc5DYOJSqGWLSIVMxeieNtvDQ7OqOBtPKmrw5qa1MLdVYN4BBPb+CXKtQ/kEx
YxBb6R36qZpF2zjQtN27+pZN3v2EG+IA3b5CLvjtpkjY6WMRWFFFg0R4nFuieDASdBY0Y2ufD1uj
FuZxlvH+4sm59qJwqyLKtshIHjbzFJOX50H3nrSquLbUSvBoLLJM4g8a/Xuy3Q4z3bIbzV+l3TKf
LIBHyEasxjLO1l2+0PPXerSW4TSY/PLcw4MNeF7naYIuzGiyknrpHNEOrEeCCzE/ys0B/rzDljEW
JuSDKovewhEZlPeHozhO3pTlYNCvZYJN2hZiYUromzwjAWKYyFMj11NYGhBh34IDxQj+ow+UiF41
lOXjJCJ0iXo0dmY/xphclU6tmbuDEnpxKn1tRMIc6ZSmbb6sNpbn0ZVsOHveA0Ob+RJqSX6Q/Uy9
n9XZ3tfZZh3oRULHyr+UXY2w/nFVPNgcx/xFpZ2GhjrjCnn1SkL6JRuBMDIgCcpGfuS/jCqm2Cj7
Ykj735lLX3kDdmAp3ymk1S/ftaAEmS3L8jCaFyw6dQmbyu7QhXexncwYVnZn4/A+5kfPoe+7du0k
5ywDKYuw70D3/5LqiyKrdNbsjVvV2oMMuVAt4iLoPX1p2mKeVSmOBXqghB3dxDaHsvk2yk7ZahOG
wVX/OMDxhooIZeVlmQxIlobeYd0ge9+0vMUJfnZrGbBvk4RsWSLLUSw6NSM9ytqmuq3kpdO3R/O2
UAy14t617srV6y/m5VRDfTk6u1QWZkoNWzRmq3eukMQadwA55fRo5+5iqr/0+EMcMGwYglwAE1dp
JmZmHcfMAmpyp7Mt264UcEiPch1RzoPkGtAaGLsRL1uS632XCy2mqkPvECNpLCI17AYL/Q6CRy/9
T5zxjzXAp/79xpwvgwrRxeeHk5hfn1fBhUmXvqDd7ywWoI+Yeu50epoE8Map6KhSyebC7a4MkHvz
x3t6TjkFg1fBBKaZzD3rHbAZuzfhI6ER9RoiUIjW2gfrDUtaJpe6pSZ94BVL4mIghRWbvBp680ic
R5AVuskouAqpDHokhWJb6CBcIoK/3TGmC8WmBOLOUsvN/iVuWXzReWE76Lt/mM07crUY+CXUAaF5
YsH0jNukIqFW0X7cgItCXBBhdwrfrvVslz7tIK+d7teP8iIzeJsnl1nbTFW0yEoXXCUQhroKurGw
N2FXnCMuA14v3GdZ1BOEUHE7iFF5ySPH3YkfQNIkQ96MbENPc2G8EcCF2bBmJeVHMpco9mASoYBg
/5Qoffwz2wzfiHx+TiBy3Q4IxEBc5GWN1yVYsa976UJMyJTRyjxTPqQt0wJ+iZj6C3C1xXFhVb5p
COlRBa8ewyuUcyNd+8rJz6hbMH4reGpeZiB5pQczLsw+28iv+wkjlEHFJYKpIHc5EG1Ov+xMfIw9
jleSgzXPoQAE84BppObtGHleSTZ6GZSOIdtLylX1wPp9fkFDI8xYmBgCtoAOwcWLP4Vsz+8/+kW7
GO8NtH/Kn544xzLStOlkN/jlPyYlspXFMN5NMjoejNBghfmK3VnAidRy5AUobVb1EyfcEraC6d+1
k6wmmdVEQv+AF9Niu9mMOBNSj2p6eDlmzvJ+tTH68auu7+Tkp6rOA9Fy/NEddk1wyv0ylcExrHfz
4chD6V4KWUrvCC/dr+Exnbkq1xLLlF4J67sw51SmCD1YOS16yqpM4dRQtV19FyeN0t+Le92XOHLO
tETXbSWXvkT4pNpM5g1GnFek1ae4V+DjXlwPKNU6ThOinpwBdtCr/6Oq+QMnRQWUjVB7P0ummenH
Tc4pHYIZF348xYTLT8zBOdxc0DVoh5e9X3WCm1UmZVVErtB00vX2QqMbfta0Z5j4amby41zGdi9U
lm2sfgQQ+JdD34KM9udxc81X5Zi2cz/uFm0LCWz2v8BE6hXMOBd+ABIPLmZtJ8bRmHpLmin0MZRj
rYOdo65/emTblpLp0KsjNdN+9BeA2Op5j05ON/LqhZOH7YTFCPhAq+Q6QSfRgJgFigWtCVWUl/8T
CdGV9sLKCJL96TKOd+Z8Rwql+QDqrnyj4kFLORPcX7J0BOjAhXxalR14Dgn0WdPoIo8KQBVkP8i1
ze8PiL0g8tByysHp+FljEAZAf/fURjPLK7uE3mYbkgytcvT5n+a4z/HW0qcoEJkrMZN/HulrFemH
nmA9b9f/oFTL8jaLqUBMwtvHBZZaGAZnsL0ycOYRyae0mW/NBj2YTzE2tW7J8umIKr1BwmajR7pP
hPDqPH3lXEF2mi51ayOB8JTS5l+sOalAyZzrTJgpydLsX+j6zZ56icChQx7MfMjvlGmFfKfTk+gx
3TO2aQT508Fg2j2XjaTGFAmkz/3LXUQsXK3OF+B7s4o+1oj8MSdT30l/GQUWA7t2xZGR8P8L41nN
dXUwwcFxcvNO4N402vak5YjECOfK2Wgg9U9agik7E0avbh9UMAu0YxpI0OCS6D/Gi11grKO2f9wi
mo2M4KFn81r7FdVfRozQIlaOQ6yysPZtWyKb+/d9SN1ZM5iwL2ZdFoLqBawoA/QI/YN8s/Wvnzz6
V4f/oc/iMneA5+FrfYlNPtRjrEcoJGxlXrLltFAAW7A2iRPQs9kXmSl1sJsla3EhXgML6h/c+wBB
Wny35zz67/4W+AwrvxoCXIEu4Q2e7s0IGhS2wuCz1v/Wg1bGcLOkoiDqySSSRpf+NuyFmkkT+mdB
GsR+TaGfW8nJuyFXBE1uLdtFZrOdkm4ZPXU0RuCBKVF927fQxfpxTCBicafTuFjXAdOUZoWSPeTp
4HdYubHTKBlqbUSQmiHbUvZMYUVpV8lARyj7vwBiC54uSNBm2v4Oe2eANIZ7djnF/LK99xe2fSg7
/+MQS+5eKLMxZNTeVhVsp3xeWQzaO6/6PfMqun9VZGP2ehADdLJKjxHv9h/M5pRqsZI8mndka6JE
FgiyJ9eeVrk54Xy3i0qUn/Hl4rGoymkQCm5FE8/Ter+aeuC2iCEEDXyGZOuvb9Sh3je60vugKPye
CkuyjSf9NiFy37EJ54PKLuSf7y/9w+fu9TpA5L7klIszrTwbD/lOC1eNwLOyXDKqLuX3mbW6l5zD
y5GJPiDEFGjX/LH42BGnZ2bCm9FU/B/pxAmZu/tihEGT29sMHoZd1QqTXitUSB9iGq75+MThOTmY
HDan9ZJOMjgvsKrjVb/nPClutcfC9VKypIN7ebAndjA89W7JRXR2JX0JR+rlWtejCq9yEA9/yq5r
hH+rnZZHFCjNVgOubyFzdHoxttQlIRMQef9OP6xWpHtfdhoJtS2qpaicQDtq1oCut06KBwdOK00X
cDMLHrdCor6RoOfTiaOACnr0oZxu5ca1MQc3OzFfouQ2G/KMIx2kWGoDf0HvNR8PKCNmWmsw9t8B
hjFKlkwk290jPcS4XCJ0ukfxqyUG5ZfQK0qccro8l2ZLE36re0S+YqaIOLBwwykhQ22IvcmlvzKg
HYnFEFAH6PKVZ7oVKHOhUwye/b4bUnbRiR626FSVRhJaS+wDXdG7wXzCqEwGx0TYnawoM+CzsIk9
5TbrnaEYewsVk2WLhgA73sUfeTMKUpj1wA7sdhjkQyF+R0j22DhG9yHm/HDB2S4SUeGmXJJfe9Pk
pasf4xdb5q5jOvGC+nDQbsQcY7TDTI28suWT1A1ctoepr+PUfRPP7c1dyM/wS480GTrcco5UdoSD
51TO5XvR04JwREf2lt7Roxpb9gQ/eOQ1edxjDp9ujiovDf6JHz5YvNv2wTdRSyJL+IprH+OYoYk6
22Yp8M2ojfkdXz+UPII5bFcjXAj1rZ5tRbuBOYYn/m1XWLzkA6ljqYK+mOugTOy+9Rf9YS2ABFyB
HC9HvaFfiLUXJtzOIeP+XciRHRnTYVSjCGXzQdFMLQAbqJJxu5YKCIIcq7MHVCJHZ00hNogtNpg5
HWV5SaS0CFLc7Zq4KtiersCmaC007IRjKjUufCtU4OcnzdmwFggsKErKBfvmUlnLLqZ2CgkCPVOX
OPM3z/7R3l7RwL/TvvNKnKV+7EjTF416W3OkO8HhB/Yn0UewrtDTCf7kQqitw98XkaYPccI4eDai
5rspQ24ZqPKcfkL6X8Fp67tyDCd3t+hnFa9ekygxsCUsJMKRcoV9wCFgSZS/lqoqjWyR3b2NmjIJ
JICQz5LZAnjarwE4HTAe7rxADNEl+0E9h5BLCFtykR8nJELVU98Z1HRnZ5xwMleA2uHFPR4XRQ/E
p+zpqbKBnRcWuvk2GEVDs3nsGX/yt+raY3fcZ6/SO8xhBKeJ1oyHMBs8Q6scWjUGF0ykAoGncoOA
KA4YkIktTOJThcQAE8KJJN35q4+Yh1lN9B1PDDW4cFdKax14FKU3L9fy9FZ4wFm5MOXMA3tpqMvh
kuA6bpNHBbbHSspG/0PPR7zC1cJsfH/VI5+13wmuExuGTDBUCzV8DAnDgQY/CHDdJr3rcZHrR4tg
bAAI6t0Ch3w/tjRB4WNOPF41PDICaUVZ49TqeckWD1wTlk2tMqiPTtRZ6LxO2EsCsmELw40nN+DR
0eoQz77sMKJ0ZRKXcYlKkLZAvxL01lJT3a7TkiHTdgpjLJV3F5teCuNnoqBZ7EyR8MM9QM7vVMKX
igsRejhyTy2gJeUGGbiRDxvKQUdcEQT01P0v4rQW9SE0OfByIiSpFhiiZe6yXZUf6zVlDSz0yhpC
fvLbvL41ODcwx+FmrNMG40VfBtwjpdCRJivHUrZF+lKD/U4De7t0sMdStJoSKeGYtxEUHtnE8Cqn
G4tpZ9QUX9mj1Kn92nFdb3kILN6dK7tF4h0iTuGz2VFG8p7hslGlofXTNJ4TQ9EYB3c2MbfYKHhc
J2cbCt1MC6rGnCZKJ4X9330AztD+r8NJ/WknoIa51rnbdb9QfytBRD6G1yNatYvxYzbUZIpMcc0R
p7FhW+kx9qScxKCXjmzJbrgk8XdCB4CTEuXhxtl/lrY72toBudyVyqPzcedIsPHOC9zGU2CjoSdS
FZwTWBi3zMB+YGrqkRa5JLOsBg4VZjH9VvOk1dGH4KN1ZlPhWa7hdcp7NyWo6xB39lXwYWWM4qHr
gT0LFQBuxPe9GHHuHC2vqDgvkd/n4iXlx4ulG8heoPHADUUd6nAI/XA6tirBxOwmgxTE1iOilWXF
7GrnAndpOJsRQRQljHo0A0TlxuPS+ZJIzskJyqg7+AfFyBYFYbTWy/ldSukycxDQbiHKtS4MjoAy
MGz8WkxOL02f8diB17n2mYb+IeDP/HhPyIkCyyLOot0uFWVzAmAWqhzwXrL4mh7qKDvBvC0eF0XE
VjlMu0SY90aYDabDUUHe2jVP2Ukd2GxtR7yQ5uniQUlhYA/k1ir2aUUVUkcYPQxHhgc08sjqZ53S
t03P4WXencwfWX0Ed/zPxLdMytgy7ytKv8pGdWnQv3kE6lgQnG8/KwHW6/MyoKKT3twkPF7wUx+M
tV/nKSGZD9GCCEXNuDQRj6+QU21h+5rLzBSCKTObuXihXzWh448BE0xE5LG/ObrqTt6iBwPoJ2jt
4h8DXIc2vKRqDdIeswEA1fflzdW4gHVb7P/V5XawjmwsPFWTTcDkjXSci35+thCMgMfxGbxhJoM2
BERZYv2iuY2ibFMY94D+jRSIiuZ/q/wauqWmrplWMf6gboiYbq0/FiSy4UbvrFcvQV8qHgDGwoTq
riHC7aVSl07TfJpLifVqsVm7mV2H7TlIQk79NtMO5C9n1cKB4R8+uv8jqna+Q4FUMOlrTOb0cUlh
rxitxd3r37QwkGxFLwdGZqBcx7dCmwtm4M5/SNe2VnMRU4Qjo7//sOoqWILq0l8aKSps2IGHzgg1
I7FtjWTsQyizEQQu9MfxtIN1DIQFKpE4taZAvUeJ+r96wWuvv8KgaSvBxgWMVDnss3M1bKRKVtlx
e/c+1DeQ1cnzlwVVlYZcO1tbgJsp5eP3GjGcQD+/F7+Lr4Y8UeHiXG3CVxXSzqZDHRH8viZr5NMv
8nsq/1BbcLI1kdqG+M56QWw+U3V8xwxGiIvPr4/1bP4K7NzvBDwbhY1lCymm0nkzClANG8u20/Uo
Lmer4o52P+PrL+cnWefT3Dme1k49dnwvTsG1SGOkpwvq8VQr6fTDGoCOkmjYZcKJYDPa9PqusRnP
H9meON8+CUZwHc+e9BEVjxNfJ0pp4OGy4r9TsHPoREe/eJNKXjGZfxZ8MpPI5Wz4v8yQTN4EbB3B
45UZQRQHPIqYyRWUw6DSNase6REvLkfMtXvmoWpT8CeKP5PnQ81gUY38wMrYplB3riZsVvt0ew/v
XtO0MzV5R+fVU8hOpaR3rZn2KZDIIxAKzRK9JrH33uKwE59+CakQC6NazcEQAXeF6vFdEaF1Htoc
jnFwiIN8Qj4bjGY4Lnztpy8Xur3L5FrGtkqNNQVk8fuSBS7mheObmf7PD//zjG2nrNKxuNfmRfKD
+lbQna4f6reCLAujoNYc9Jp3MCnEYHuWzq0zI3ixVDYniJwj9ylGUYGoiYBaTvDxZMRlija80HaE
vxSGERiSDOdgsdHjAbaltCQwsrCtC3rXn7888aWpYmhhbgrnxTSd/mu6ZAa+SflHMPYUMvWiF+aA
vtRP+SiWw4loVzMuO/3Th+4zMR4Spv8l4uYg0Bn373uORCaD6ZgF/lA10VEIIoIBi1UCw9QVCkZo
4dxhNyvdDQXnUOarMYFjN9nWQa5jCvwI4wpLJzc/FItwmxKCG0s2247RJerQl81hA+gq6m0WQd3a
oFcbNVuO93+aKqu3i+Ph+2xOVbPHo1iK8dng+wQ6APEO3mxPK/ELqgxvB27c/bqGu2LfXixUzna2
2FzjPth53+NhSrCHDAf2VcZNUT3i6zIXMXp8v7Ib4gq6vDKJTbS2axyNFwxEGAO7cRqQ0937x1jr
T8JcJbwnc3Dy3T5lKVKi/NNnAPbj4ULjzJ/vQuk0coyaY4FLuhZqVJ2qEnbdKLQ6fjXLXDsQzb9b
knVFSr7KL7IUB6Ey9F7xMA01u6CoHJCh5zusGTvNDio1CZHFoqDVjbyJqr7J7ZqG9WES2R+WmNUs
nrCipe6eTTVTYN6mFaqExl/kYW7gOU/uq+0frJ52wx+sRuI9zkoGAsjyk6PmoBtrc99s5ByJKBHH
PXSJpXGOYy6De7t8SefbDKzSDQklZe8a5bquOr72U6EcMzjaIL568eFN2imZmtZzMN4iZNgE1dUg
vz+UvkrGdUWRcf4d9Um80AZRu24mlFqRR0VPQrhWxpF6JbBF5UdBBqB7CPeBERU8SphLhsTutKNr
N271pv39wC7VQPbtTBqHgThIXCLKNUlBXdi0XdRngqD5+RBlJriHGT2o1thU1Fu64MbofMIHCM3D
hgS3wNi8wHCdZR8ozHlCvP3VyM4cI/0/BZe51AYy1cT8REmhQ0S37MwyLztmlm9h+Vw2qL9tvfvl
gJX/SbOo1u93BcwLSswebjOY5CFFMV36myOMnpsoqo7JvpvuJIFZe2dEWy/2fs3D45PeoGDL6jlg
dwIsz4dZbPgn9KUyef1Itp2ssXKQbsD42qnYsFIIEwP5GdaIwZ2SwcFf3HfoD/hCBX//FPzjMYPg
ggw+0RFvxEqHQpWk9d4wfCE98dZsiA2P83aIeHVXzSxvEGH1dQnNruMdyFoNk1NQ7ZEhXIs1QUZV
gxEGiSXj4rQi2vyINlmq+gJrtIx6FXCicnta1YdMH8MXrKc1refJSO5KpgcYWFiJIUby5v2quhlq
EQWJyA7mNWQLFurKV8RSwHN5WXW9J9WE7F4+ujqgGan3XrIEBknqBbfrTmIB9D3XaPK5mTfC6VMP
Ij5XiXc2c5HR8egKddm3OSzU2cIXDivoyl6hO5iaYh6HHDvrWk+LkC4XDbD+FPySOv9d9H3KfYZV
5wShSbNINfoVgSCmKmzNU19ycDR/h+gqOmbP5mn+rZYEsPLCiRTnXjNPyIXDCD+8FVb3oFvsEtvD
UMZAUM1pbKvuj2bbpgQ06j8IB7F8PD0eUsDK1hNUFfa5IUDJ4G9sHPKC2LyYPCfRvbcOLkQpG1Qb
RYUVQND9G2VfuDlDuqVrdxVZwYagwr/bzEQve88xWUzkgMtQHUmUjIC987MHJcdWsn0EZ431gl4O
yxFcjD7tvd1fPYxFpDcLh1Uq01HKokXMu3JehH1rFugIB0pY602oQA57zJwD9S0KggGuV/7jjy5J
Qzoi4yuV8varKxPd6p7B1k0D7umfkEoZDUdUPeqWJYB0/suf7PGvNrBvY2T/wkGpkkN2rb+jhAuZ
/QXZXUSwxnWhqpKeoyYABOiOAmzGLEor4ol7n4m7CceYZHDjdoI2+OngS+2f6vZbkHwH303rdM0c
OBcHBA0msLpR5r3HQSbvmp9yT4uGtGjZwcQw3eKrGXsagvZc8USTlf03lpYPt/ulkS2abMC5CFFv
cZsItE/jPCcHUkfMLzDJkDorUat7IECIFH385m7hgh1QQze2iEHmWoWgQ9aGZvomrFL0hUFsqxJL
GUqnaSaOCP02pBUrDFxdFi9tCGX0fQ2JOrAIUiTL4xg5tkQ/qVfggiB2yix6TZvi2ZnXzgPZI2yJ
w5+2Nfm/ZNIyDd6ZsaFcMOOcHaN6xQi8/7mPjkSfMuO4EvzVzmLpPJTSs7JdsvBWeljsariEy+jc
SQgfVIltrvykwBtRkfbKh+qd8TmJGWMhg+Qn70s1ezwgoQOoHASV94hlWPu//F/HWX0ybzm/7hHm
IuizrU7UmCa/o+ibTyDy1zkdpAMvPOakE8M3Dc1CSNwtT0frDZbJsdP/Wu1m4TM/GvIU9s3He2WV
6y5ns3VPEXhxj1OpfvlmNTUoev6lCdI/aZmun/rAFQmSUk7OL6yz48xDtNz1499gAvbUC5FpfOl8
2yfHm9WXoE1GaD4NQbNT9HZrZRb/SjzGReQpCcWodpCu2RslbHZ0bez1/FP/aNF2jpub68hggKBF
VnL9iLXeNDxvuMMAU3s7ewjbnwNWWEmi0cW+tiNnMP+fudQ9CqJIvwcmx9NR1sswp9ePtr3CleRW
E8RXeEqqW5zZgrbJdBSWY8zVw2osQ1YoRLG4QdJlsGPJrp5nsINVYD7KpszXaQ6UJir3vN6Yz+L2
vjq7gCL9X9CH+aLEfDyKXRFU0OP2/1+gjGRY3JfM6oQPMRV+eTT350OQq46kRtAScptM/dACcTNo
eqnkhDi7baxy9mjnGV361Da15OEKpNrb1B7+pxWH2HlFsxadArJ03gD3BgCJMHcv+hVbKq2ADZY1
h6blqERdPsnRsB09Wbcn5zM73CJEY9RaYpqa0+np296HuQDQCOj62QuhKi8bF6uN8GIBxU4ZKZ5y
jtQLEvirfJCxvFs5pJF0rIlqMAa6FsRecDVfIiQ2PGkAUJ3O0/4FKT4xKylF8ZWk2jUiC4ckJ2op
nsPXP1irAefKIjtQYKq/ahT/UMHCSLxiw545O4hqRYZ7AOe2hE/x5J3KIqzdlTYWe4aEiE0hahAM
giqMWZdgJvJbdtSDMk9iLm1BeHKLbMPO3Qrno4EuYgbBTxXyjq48GnD+So+bJDCXCz4VPeHlkA9S
kaslSLdjj9UfmbwOUtwuwTcFym15JRaMqtZ/at2j81TDKtaKdUxAJch0hm43OS4LVgZ1w4siPpMo
S2JF26RI4R/w+QBX+zCd4eL2R+cn4S2UjbUASOMS2A5V7RRe0QGdCIjaBUCwrAHnsBnRrtAGON1v
Nohobjzz3utTMTQAcEnXrb/iaKoY2aU4z+MseAqkS5PnmrurxCFOPhfnGJghnGXQFrh+ppeWwSj4
g39eCQRPFrkLOh/81mYoHkMBNa4HLkMD+P+Ra9/FD3UNx3suIAUXcjnzWqFqXw74pTbtLN/GQ8Bc
wB68uXrNdZRuh+xvH48KUzO+me75iHb5pMC4LOnBgYmcw/RAuaQiyCGtl6whaYQcxn3ddwcvWvB4
PVUvHVmDE9pNG2mqrsmDnKpm+molDCTvtE4x5BMXvJAtddzpyTrM5RqJpCNdlBZj/bR0sM8p1Wu0
V2sordck86IWFJBp1ixCJC2jPIS4a/YHwmxoqVjuCBZmLeS8WxLAVvpfeB5mvG/5EFCXP7jSPinw
15qNUy70JuqjYH90ReA2PXRga888MUDIEETcd0HSTbT04n5pgnjuUAytyEqorL2rHB0ziCGGiJS1
am56a7VjGP2DX1Nk9aA1I96NvlOJYPfW2jMBaMbxRgZ6hQ7FgWh4CYGrNczrmEwYajxD5PtRTGi7
uvMOpMmsgK03ckJEMw/e4OiteUzo2bsjuZnvdf/ipwfajhelAfsGvLJgcuZP7M51UKtF/wcIu2Ao
AJxQEGc37OhFOdeeg0ULA5BgY92SO8IDvLxwiA9akeEuqaGgxLpYm2TXNIeIbGldK9IgYslsSkpJ
N/t1heQ56H4wCG4JOkP+aFTeqqxPc7X//+s/E6505Z4ACZ/nJAqK10AMUpCd3jvQTQouqs6iE1HE
sgOOQEJFukDXE1Bc0t80Bbi3B3jAy7jszKGwGJHS8gKA6xGVerHhjjqq36/uTrkX17kd1LrPV8d7
uAtamY2AxJys1QFk1+1XCsxxjQrnXfrq+pyya3WBsbXH0etC/k/C7xKAgBeZFVhKIK3r9RODNAYG
+PBvpb1TIBdgz4ua7WzFGGFBpLv3JkJF66gKOBWXjo1rRihHvuWAca87m/QBzbPSXYlSOi9vk6BA
4BFIglBB0aRo3Togdh/fCy1l9u5j3HuvxPdM5YCGm1N7rOFbDPpKgkj97kQJWUbMohTgSenZ/5Ik
hSEHB9t/8DmSmtkdGjMIWuEgkp1dPQ+an7gsBMxd7SShycGx866XDuAFhms9IeObqygy/OQtxRXy
frRFq2lovkYB9pRK6hyrUKsSWtY6tmt73+3r5iJYPansqzCCjuMdn5OHZFOiib1tQKEOWjTc35oA
2YYELPf36QPIR8DnxSnH9COGaG7Swa7MIH6uuckOCUZglXmp33bEbSzlpgSMfBpS0XNBpS8A9tFG
Curp8SsAkeytgSlkMW6FvT1ShhHCcOb2Yy+ZsnFp40C+WIcn/fMJLTTX3HNFWadL3J1XfcsMJY28
gm8skPioE4zgwTjdKjfviG3rK7YFdgtjWR+9DxedF/hEmPeu5NDB+c9liXCfnn6oHh0LBsPzEnFq
28f7z+S/S+bfywuvrmLHlunXd1TKHZWocbWRvKXh6B7W7QplVBClYQ2Kn5vF+GO/D60ihN0X23EU
ZYQS8hPLHnBqZSW00ZOEcWnmZCCSS7WfcZ3Obiad7HmaqIOKFZfB7doH0aA7IfTqgBHGVt27gps7
psbkPF24TnXsuXQ8P3TN78T9sp1KgMWz/izkhn/Gf1CY6Kuxc94V43jH03QDrVvWiYwgw/V64iN3
5PJEI1XxfxurbwNnoNuMkCSRSNGqhT2zHef6LJ2Sqg1IK8gJi4va4CPcLUr9MkButx9JaH3Z0XVs
2SpHebrhvBcF9Dw2OnlAFPR5CaX2F5eN0JIvkOV4WMcXObOkxz1bYedEP/IS2RkvRMeTd9xT0T71
2fUzkk3zic3MH54cyFV+SzlCUKpVsVjTj0rgLYq8/D2PBhQRk94PPIl1EeB7NFgg/i8wllrcR7Hd
PxmxlDuDGfIX9XJyoGO2WpqDOVDPxMJVBLfY15HUkvmlWorILTKCqDa3iLe2FzedctBqRuL1UCEe
XnaS7b20A+/3HlO2rIUyfzJs4UG6rE1uakk0xmaK2y4Py7GrY4S6WRkazL6sI+MMn0rNyl2SARwd
9uTSaKf9tgyqgkOlzdJ7QPEBUbnL3q8F5TfZnKyA+H773dR7eZSBi9dr96UA9MyzIPZ3p59MMgCb
Ci39wxyA8ScKGovwDmxmu5S0FR6I2vSzI485/MBOzgaHk9NTJ/IYOLB6+SwrFGgzEsFiB3gC3Si7
LbPDs/Rj6FuDvYyM7l6rtMi5tPh50j95tJAwRPj1NPdr6M9Zonuec/kY269EtpatJ2+4tTuQZ6Qt
QCE31CdAglutTtd7WDeItrmiUvr0LaDtF/Aaod+ix7fyx3e/B2A/13tkXWUINlaee+ZViEzTHu1W
3sNQUBFbRzczSp8eA7hAID3BBCdxXakZG/nVcb7sMVC9IvXXG13BQXcBTwqxl+rfp1MoAxB+iCGz
UGxi6GTZmjwq8NE1dJKCcY/HMEtqb7LVt3pR3jSKeZIbJpM2XRm+wBB7ZGbeGbf46lE+HhF6/0Yo
F8jz4TCBuMUqN9InHRtCc2BCWd6Wx7/HN77neHit/CMZzaSBmeHqTF3Xy18ZmPIAhn3QX6GdXnf4
BuEQ4RT6fnfl1JTC21Vsn3Fc6942ueAKhXisi2bpLHAUol1JcrX17SRTv7PeuU8Zk1gDqQ7OUM+S
Vh9k9SUW6alBoT1+fWYOLCyjmL3OUobNU8RvPi4HIe1CDopnTugljx0tBRIwvOM9rMNTY3KeAXdT
phTRCT5mfQOd3AkFHYNbAFodAm+JqrsV3P49CvN+tEk+mboPd3QfqxoNyEb5WRSrPrt0t2FVRIx8
LxyG1nC6CuXZU/AjduBr3WnrwJsigjUdc2ENXq6MFE7KWwPbqZdy+CixR8tsvb7DfHgHq+sjF9lH
gf7Trryi3pgsfBJlWMfIMjCnpG33txbK2MlhnDlG1D4+quKUjuw6DST/T8x+HLvOZ15OntlmyGL5
xR+yUGBLOnnolkM6bssf0uLnZuj1lgkz84LWcFDAzjxjezbEUvKx5xmYIChWKH0ODwTW9bDnUnKs
i4YQZp9PjKLBJFN7R61rO7OVwQXGhLsqOgEgARuvbBUUzze91OS3H/ihXumpWY/oIM0kjY49skU0
AhHgGAb+QJSPv1Zhn4R+ltVba0aw+63EOVvx6oBUezm4FlDOYem9p+l+3yjCvTRglAcqUFWif9Cs
2pLMiInuWuJdNLnfgj3ddfxaflLSnqzl2sLZqXBPkyLiVj7zVPVUkE1+cSLlYLGDLIoysIP8BkQh
EpCPa/PuA8LeJli5SN8dDl9eJIQBipGBcRjs69AhPSHWAfIbRdO2CRdns5DzsZj0ZE1bIbjxkXti
EJ+tJ9bY37J49Ykb3REyaHbM2hqxHo+ApKrbbLGtekzwNIVyeQzJ+G1uyPXep+CrPyJ37yo4S88z
oKu+FFX2Xp0J2+QLQ4+sLp744TUtmp9GdBM3oiibzfK7dYNccz5qUZfOWlBBdsTDfqG1YPjNLlBg
1BPAeX1i33B15lEGrqHFwoKwTJ5EECRxcja+2X9vl7Mt3QzYfxkPMMBedpmOk1cRjCZyxenQxhcm
kBIqD39U7b4cGNrG/IviPycsPcilshN57zVP4/K61d7K3qbcyiuyucouP9reK7YKR+4T+cvLsd9U
NZmyMLU9DySxNTk4UZKssKlTCGrgeYydOg7E7CWhFdXmi+B71BKsZMKux8dQqrzQEXKje+caaJQb
cFvSGbDL8OTbYOWNv0F+4PCpB9ofJJb6ntzuI4oCH5DK42R/5D9LeVlVXSQd2mqDf9KhhK/Z1ruy
Czd6idjQnrgwFGvi75THPXPNeBD/LbBSifH8kO2eTba49tGlspyws7zWJIzKSi48nkz0DsF7a+AH
fbPM991z5W8AfbSXWYzd+rX2EnKwkYtZCM+hQYSWX16TVCZxImXzJ5DxvXNEtpM5qkC0/EkEPc1Y
Fvro/lYSIG7NzVypbpF0dQcQ9/5NXSILaSHc3vmlOdjzA6EPJ1T6hXVcz1qa/ETNMFhAPE7zqXrC
FbDwdstxRgLIJXzBthTsd4fC8BTZEKQoMVQG2OrB2DG51fakEeAQACI/WHmMcjyJulJMe40wgMYe
ny4U2jud+39/oYeaqxfg+hUi243PpoKYDbQx8b44lhyOG6q7X5cH6z5n+MQSZhX2tk9WnJAOacN5
y5Pl2ZjS0eeYHACY+jk/C/4YycODc0HAgpSbJfzBr7JHMo3NxbBKKcP5nXY8tC87+z105CZ+HNu1
b/SntFLqcSSlrx2u3qGNmncNaSVlR+HcLq9ZCZb51AhAfCkVTlgtX03UqxNR0OpiXrIex2R+VutK
o5SpOMtt+EXCjypFxbTd6Vx+twiSsF1xmOo/khpir3FdJ+oXB/Rxn4NbO8UM4HCHiu06dPzfKtOb
rS0ehQZVI1+AypodcpzXG6lIeOQSOXRpWLRUZdWAqAuYvRKxR451UnA6frYUeg/aHLFzI6P3oNVN
M1mu6Bhw8762R5PbCmLQLwUZh1QcsJ/qEwHXIjOZLqzEAy1Wlz5pBpEnV+XKKxT/2h9lbxGycg7p
x2qXjgmdEhddk07jdp/vbpV49Z6HC6zFZyMWdU+W9FT5xPbSHlliTAv4lE0OQSE6Y1EGg/HYBBrS
fa74lRMJsA7Lq+PzObjK8biaREbeSCLfkcihd5V5KJAaBEBzUsHtQWImo9MS4IMIsjZr1d5AsIq0
MHcVCwrUGF23uSNcOy101pqgIZOvGP+FzDWwCRzCqfX+FamvhewsjF1g7hP23nfAF6yCLjxe4kvn
SyxnWkumnRIEPWZ9QH4BABJJcra3Scj/5vA4TS78ZywFhtq5K5cfmLqdMrYv73TOPTwstbYs55L0
ZwaoIUxApjHa0km+ojeN1MSSKBQ5clfUlvtgCCrzHr16liaeOsq7EoffDYUmI30zkUPmSQ9W+9Eu
+E57bzNk0nS6orshz79vQK8Yys9alPqRRNVKiidbOH0+Dkrz1srM3Ygj2QE134NNYrXT1PXejZmh
PKSpoG30C+rFOqGHurp7OhOzP+7pH641du4l9hg4wGFsmzJwRIioXMR+B4PA9ONYaopsfph3aKLb
Fgu0ZFLKdZQoCNyLR8fAtvqYq7eADzoE3KFmt5LPWhiRAV8e046HIhVz07wsYGBosuYyVbLoKOKp
cOU3I9JvdDwuZogt96HKjJ3/uGyinGkENsWm4a1sTwubjK05vhFacaqB/Aez9fNbLJNScLXa9nt3
Hnd5THbAPj1dRrqe8YSUFUN+z8WiMzonAbOLoTTOYSnKnAupFcFktkqbTCjg09E3dihmzyDnro34
KXEPFSLVnYx5xVqwKWHmKcsw1XG+vuQv7f3W2r5qMtD86d77LZFVS4B75d4CxHlFXTUmv6PccJ3e
XxbFfICyDaoLKbsa0nfQAS7PkWtoPUc1H20Huda2LaiUKXMTv/FGfmrbJQkPaGh9Kha17JEd8p4B
kszYliuehmC+9V+J18a0lgwQr0N2993wNILnke2E2FEfXN1svrGPTwLNc2iCvmeMw9g/wfA+cRJG
oUQUO5tCusMbw+IwNExtzb6CWzEXhUmaHPeNzyjAYR/ZEA9dgKu0t5pUoWIjFQkCWGsFPsQkORRF
fP9qtVcLK4To6BNsniszEn6ICcIjJU0UUmuM2KIhfUESwMMY1n1p+PA6T+4FsSySMeo0oHFou0AO
LdtkibOqeR2fTyohSeUnt6Nq7nOV/1k/s/JKBtP/V8yZGtEqTVS5eUgb9yNtpwXzIy/gc72pd6KM
kEzvv878HkFnJEdVKx2baymhRlOhdrvVP49wtk85ztvUaouJ/ot3mAMetyAlP+HT0pz1F+zwYwWP
0YdplP7/UHlZoXAxF6AZ/P6TDhyxipLtJ4TTORdiseBvCeSg0Dz5wPp8S5iZmuG3SJpxZ0pvrkPp
lIQpvvi6Yzxe8bhSxDPJuxJ6WUgKZn/Fy9ea8edQqJe1uyzefytYYjO0SKn0Ir2LT/YGv9kbN6K1
oi026E/viElBBVLagoZQHi/FFDU5QRas1ODI4BoFLNq/H/vVlrId3YkJryPLjv60z6gUYYUGiMoL
U4FeL/JWaPM9suTX9V3TU8Hw2tgpkJH0vwNm6OB5pb/yYQJT1e6p3h64uUzzuw0hGtYEfeLA4XW4
PyQLRahaMJ5bQ1HTIsKIZcG12+9lcbPoNT1xaMwis9gc1fw8nOSn7/MIX6ky588YdHC55AAybEmT
dNiqe6vmLWopnNyCWJES6gY56C0TYRk6kVRNEyMduuaMZA68b+d3AMvm+EgCutCE+l9UPuWsWTuM
OhabPFBYJef+RaazVdMDNd5/szVLZmIaRgNTvduhphIAEILnk7Kr87oOjKoCyZnI2uRDDl9U1WJp
EYDanB80+21rkE1BDBjSMAtZ/J1tcR/8CSOIyyPrTC0AoD6hknGYUXqWlazJiOaJjax1MJNA+uEk
mXWsnz9kINBKZHgGz4mArmLThpQuIgR/ARCcszDqfgAEfvoSNc43A8rcwE3lXnBNvglJWVPxDICW
T/I48k5Kj2MofzY0Wxq2RKIUhXX5aHqXdGtV2/ybKYFDLfopXIdLR6rmN2U7TIpvS/ydSRjtuuh3
XC2qagk2/kyqoAerYcjHwan+70pLLzMMGNEQ0BBUMctc2fUidA66n/bOZqEB+Z38GZlPIfEO/eOt
kA+CmMjDlstD0iI5NhPK5yGihD6WS5oTwf9Gasyv8ewbpCOJ+rTWJniE04VxiiZEXCwskgXyc8m2
l+aHBl+ujca0zrmA3NlCOPiHQgSv81gY5ru8aSkXOiiZe3EAkQkt2WrM6NTrUbeJyIQYJ/CJWYvF
YaSytpUBphTwOpFATh/bXWAQas9iSnrn6PKLSkx92SZCHw6Nrnv4KEEQS2c4SoicMM5Im9sOjq2s
5ko+OH0X9kSSIcWfe20Lh8Lkrw1/lCl7ef6Fnz0txtoBorS8bTfQmOJoA0GZRuIsAtfXVKZU0JLi
UelJVfie5veyt2v+LcRrp9ifdOpbuaAO7X3demKfP9/qmYGFfS6sKLQ9yySRpd0s6H8ccR0lvsl9
vKDJPtfC/Zrf9NU0TJbWsTyzb/ZbXncBPyH55yoU1NDdUGCdyvJpIPjk5lu2XUwlidkCvUBXbH3+
19/dRN058kfO0QSNYh8bt2tbxsxds/KnAWoLu/UysNPTvDkKXAUgWNUhPuYDZiyhjmrCEzJBBpeO
odGYCxX8CxL92blxJQmLQCqhLhtXBIVTsDxLhqGW9shPj68KPfNUxL6FykDY67GEQW7KzD/sEu3I
NohBMtPGRNibq1tkF8VGgBrzwI/Q70hKfe1/G5FJSkA8QWeWCUOOkHmrbNWNariLvShi2TmcRoiT
gcZW4645MW5aLxEu9L8ZxUo+AIgjTRAe5KQQjFfdyUbpWXdQFy06lOiVMC6D3dY/MszbxPz1Mffs
0Dd5j4scEn5YsS0N2oP6anKofHD4kRK7fbuzdBZV/fiVv5HZc2iqvlhOkDEJ/aKJc4FkhwGpxy6c
CEnGOCSl+t87r8DYmRcqIb1s7qiF3f4obuWAFKR4x0nPRNZd7ivtK+2mX3jYIJM9uwdG04gChCMg
08uMZMGljUxLfd4w5+MmY3I9Serkzzb4/4Yuvxif/ywnfhABWGQOx49DlJgWTT2OKmaVEWEdk/3x
ZSicIZCj6KWY7RR2bBVSJ5D86fdbxWS68pwDwSZ7tLPWwaCDz64zfabinWEpC/BuMn7vnd4h6KT0
+hDBjJSIM9QCNGIzc5qBJp8Mwap6Ipc8xkUQTyiXfHFtFWGaXhpd495R5VUL02KgQ2nGDfg0HvGg
VJWwjFQZZls6iVJpuYPmU1Fg6nUA0pOUmO0agK/65qxL6oonaN7XhIq8jVV3ojwuGDYXi2qp67rW
cnNUJaOgluY3OeML4eIAMrvwhNxk6qbLVuHY90WFNqXoSnTpef0v84gkHK5k+sEnZSvJ9cNtSb+s
1JBRR9RT1yuLNyrrWKLXS9YgZo2JQHFFI/n6gTcPziS6CVN9PZ9dWlGlz2xqnwclp9dB9Dvs+XvN
1kKlkH23rII7S6Km0tPHBAoZmMUJWoBd8HiTjuOGpGMGcLmmwEnCbDc689sOHgwjraACrax0U3BE
iYsNj54Q4AE1a570nKQKUZeM7BvJ08KIs2hFm9QNOibltjSk5KUYkQMqrBd9sM1wvm+nlsL3jyPS
8wJ++XVWkYyDiDX7UCXcXzfxtXmfpx2ivIQpWXBnTSiMnmXzjq+/7sPz9Jor5hcwVaUi7jCrPGbK
E0sNOyWJ9wrMjv13z090R+ht/xQ45ej9wz+FpZ4VdffFm3KY21dA53X/jCZndRGS7uI7YSDvRSCl
KbN1LhxKlQRDSGq1Gw7UvSq0elAOyhm07d+A/NCEM6Hw92JVj+YEfQqNfGExkFIsCqLUxr7ae6cW
QVHDa+RJ8qx0vnBmqGR4RpJQkjfA07Xf2SNhyrD0CtM8VkVmVyfxCaamBt/Vj4S97QrO8h2KaMjq
JG99NTwpSB6t2EY0B0cahrzvEuM1E65f/Aj8WYv7hCwIAc4a4uzZWMIHf+OycAJ5093jRhqikZX2
q7pzVNBE3n+9px0xQsK9HQZh4bzHdsSkM+phnNNo4akVKya7U8fPF3Co95OLyCMZfcEhr2yIKZH7
zL8f/DPuV3iHRO7yROgc3j2WE7Ht4blA6AOHewD/+Xh9AJnz+iGj2gHp+jnEfaFKXBAQRmm0V/ph
J1sTn8tAISW2dj17717ztkl+e6OGv0w4h3GncyDHzier8XfwJYEfFoD81eNhu8f/5Lx+TulDism5
mH2GHIUXzUXSwDtvTzNBZkEwHIeB6hmIDwhpt72/OUjC/Gvh55IRG/MFjTNs23S65wzj69sWmNjJ
x3xMI6HI1ZMGifp9Bjfe+4yYZyA0LLcV5YBj5LjT+eMWuoX+RJs4COw2qrJTtv/CoOs5O8fgaxQQ
lIf1kAaw40RNYPWEYb4wOu1ig+s4kzjuz7fQjtUsrgXaH5FMm5OaLugykIBWVu97fN0adBBRd9AQ
sWYgQuaP3kXqOEv7JDfqOiqlgPrX839X2cuTtUAzkzVB7Ew+yb30SDfSzbh9IiiOuC9CSEcNb1NM
lC1gOLJWhEB0daoBcOG61bEZORyI39nKVkFiGCdRLFR+OpWxt+AK/l7TdTeZBkh8cWiedDBWhSQN
BehYJJnjaBNU0H2awqgF24kwmVJ4aynEDDO4ZTQ+Nk4R/aOd864YoSjmXs60sJEq7lBzeRNi25Uc
x9i+s2TlzJODd3L0xbclyVF9Xu4Bi1o9lrrQZbQpdqJ6YRxkUsre+JxFpchorbS96OVoJPjJK4H2
pidLkUZtnbmVBQC/mzto5CCaNVjamxIoZDJNnRmshcLLa8vJRR8DfTykiDJr1S+hJxL1G+boHox+
v/WEyRYLLt7FC4DFCXWonmKKJjdQpAq2iF1LgHFTuEdoLF9vpfMVdwRippQK4Ere9SgaUbKoKoC6
UAdrukl/eFRo/RXxMrxieqPyeiiYThuRja1iYYj5hyJJrBqnrq53FvX005EJSJUoBeGxwmiahul2
PbXfFnng0XP05vo/wq8AK0G+axdWNgXH8ix7Nuom1/gzi3v7O/UXijzReI4r3aVp05rnNWfmVokP
HXv3eHC4CXB0HsiMMpVCAJNRAdd1hRzadLCBS9yN9dfpRCyuu8QGgcC0K9o2SrDIwmZ++6moF0fu
PdolYPgHUv2SEzioCUmIwR6kz7oXIWVbKot799tx3kK+2md8ExpKcSQbpca8LBCXDf+ogW9bpYv1
TwYIdw5HNRR563TNu7CP+FHjymmpjYWYEDRwoIgcgDXsy7lUKhtDWqTCJPZm064RrZq3f3kg+wA1
yQHhT+w5ZRs8o3iKbCVGCsq98mn1rXmXCWn7+BwZaKLACFCOoMf8ZKNRi/4b5Ou0o7ANpupbS4+1
Yj2bEdLbeCro8vMAE1xCNbe9R129XqvZAPmKhJmVYOtANd2tb84aBa1iTw6JPVH6X9BVHi+grJmo
28kAqXtz8QAl8d7/acR9MlL4fhA6CmsjdtjvLxjWvuCiqyDoGHS8UTuM6l8dwXfg8ki/Iblik41E
GJN699xWtYhzza81Mu5SwdajI8uok7ydSNWVIp0TR14tIQp+D/kLQHFgLpVV+23P8/wXXC2jhVrT
3GmHQGgdtf4wssQYWapA3W4mEEJ2kAFLlhpA53v59GbTCySehILZx/jU7Cm7pn8VstSq5fN1nRA4
Z0Fm7hoxfwVE+e8H0lqaNR4eoZkq4V/0FzWqmK8ZdZ2uY9Eg0Uvpw6Ov9Q1JCkMl4a0gGRcnn0qM
yu3ist+qfT+6L5N+8xcybmIs9CK1+lnu+E1J4DoETgwk7E+dvfKWFKznxQxXVs8aO2RqIZQgx0Ot
LU+/6O04f6/MLaMrYiHA/VyMXNfDew/e/AH/QP+/KRs8MpJpScA9C1kNWD1UbyHCeOd/FBrC0SII
uhP0uo0PBNEY5X8E3qx5G688Qh4DoIKHrvhT48Y1+J7piCLUi9jSpVJx5ing2nvk6UdjgjCFkvjK
Q5CfBCMtyOm2AGX1TrPMiYooMG9fVNpbtLrZg7c1gimPFM+4DsBBCmk/Y3Vrr227HxyTtWOX0mYP
cVpFNne2I7jv0QlZjTsEB9qmAOzXRHtQ3VhyzrpEmG+IdcqF4Bkqgs4pY3O1jQQDtFhqj7KDqD6E
rz9u/DGM37qS5eEYDFWTcbKnyS0mTF2jg8smFo2KJjHByH3ZxA1+xRNr1H/NYWS9lZ4YMHWZOA9z
AWaN/wTiH5dH9A7AcE9Khs0BVP5DvfsKp/1+BC4gS2pMMk7NafVt61sVTLmHGVygXRmgVdUjOB1U
/zhL6nxzQEmPzXfnEu+G0GllQnkYmdLneGU8FLxzzwXriPCef/T9r3C4ubHmA+dqP6eufuike50K
yvi46dQ34zdJ20qmrsolhR27ypjNbSDwwlldibOd6KX3AlRs6XmhRdOO/u34ac+cjlZbBT5uvBpy
tWzaiYpv1PfrqdR92MbccaqW1D2jMTPibsFXHa3aECh0K4N3ZGbUGWGYNRsOzb1XFQ+RgSvBzc9v
2h/sHOrdBwnlU+HaC5z09ABDUiGKO/rHMDt9Xt6b8G4R+LEU4ivLfBMnC9Lq45Gn2dpfsYgcgoB/
pfuKsAp3YHCyZgYJTKxfoDrIVC9RdhnMysj1ueroB5G7l44yeG1Ir7ZyhpZBtVSYe8ePlfb9gtUe
IIUbnvEe7fbgpMaj9SJYW7eaF5T4AkBzSIx48wDovqxT1OpwN/iPUpy8jwXFg7YC87qk27DlPeUd
Ptd64ESCvjbyG6x9jG58KG0vEiem+GDn3rwnZizIZwnUu/NUuOutCENks7B2uPuavIyEDytgE/fa
v6duKoQSH9DW0iVG58g+ELgX+idwlrsFeN6j66bIBKHPgaoA2srDE2j1Tu08z53zsvyh0hm1GC90
39ZcOaIBxTSF0ObMoEQchklPI69ZJ29XAkdfRNEAklnjWMfVTLfi79MI1rMmTtQK0qs8IZ1t2lw6
vE03XtbVy4+kUiDV71uRp67UOIziHtUOoA09stgPMf6k6Dz98MPKjIarsWH+0hYjveRiqnoJJPu0
683mDnDWspQ2BKc2g8OFyanEV7mPnpksDmnrJCa0wvDblnz+6eBuJD6CZsRprf+bstGZLJMlILYn
QpDm6niYpqaybZygsT4mJwM/twJLECJNwxXRjQeq9vhPcUZHKCTQvdGyClGrTqtgFdHm43qKRhun
P6quiPtxVxe5x35tu1Mdj37ZUGDDT4IQZL+ru7YdkW2ESG0ddZ9qLqjS46aGdsReE+Z8LbNt0bHa
nUj9miP2JFuRSjuk+TKmmEGdgaN6PugtmgX3yHaQNN8NEr1KL7WxrJhlzSeXhWODr/rCiE8Q9S3d
W0KtvEZlgEYt5ykQiKnq9cC+xJdJUXuAMB4gRhjWkI0y7e7Q71Lcpf5taVq1dKiEGMWda63S6xNk
nJV3y03nMzwkpDGi/DGkbRXlGtm2Ua6x+ri3vDD5IZV+9qg3AypLKXCDiklYgsVYoNylifWCVbCT
3U3fbPJWx+AikcUA9AdsCQe2t/J9nYVGrJ7yo2qcEVNBr9rjSvH9nWR5efs212jm2P4WN2smJ0z5
2K4+vI60vKSvULuZhdqhj8FmOQ0Ovh5C9qPjtOTtqpkGfN66KmJSmx2Bwr0T404KMY6mBQ6Fssvy
X+M47mK3GTcZq8n5p7srxpwq3bSO0ct2rrtSKWeALfO/nFteMC0YqS7+YjzKx550LKe0FQoNsY6g
0nB2ZSoMKGWaAmomLm3ef7hxSLI+aQLonsw7XkFr0hNa/zFPOL96rPwosdoaC6reTtfiftlc5UZv
OKn/LKsjXA3hc2ZTNpKhZRidRhocRNLsaggdNTJrdwL6+9SyeSVl8/6Qng0PCNhDuXIHU9KtCvYW
vROqcrleMKJeXaK+yE1SxjZ4g8vvKx9xS4pUuiiqRGJraxhe/WvSEjJUFK49P9h0pxPYrzm6Gor+
VJWXjaUhWLQN8IUOUwca9UhEiJ+yCAvnkC5fU1L9Do4JEQDAOL71/qEaFTp8/WbkO+OqFUkHNrrW
TsGyn5O7gVdDwL0EZ2FmCu55bQJ7z2adk6Tjyn5TZ3ICWQMBU1fpyh3PaWgXPC85KhaPTjnMZPfB
j3mYeCY9a1yDqn5tquYIOu8L/r/GHXopGTQkLzKgcOB4YnieuGCNZPyxsJcb14EcXzQex31h8oB/
wKieKUCyk2XXgLOTI1v/XejZVer2LBRjzWmVGowOLLzHxj9G6/Uhk0T3n9cm48iQ9YaQqvAtatqE
VYFcNU4nT466Zh0CTjWMxniJzyXj4FHIHPI/jpFsJvuDmxdrRDy3ymID2VA5psOJu94rz+cObI8E
3J3mrpDZqMQmx98sIq0yq5rpy/Id+sFt4iyK7fG2OaMuyXo9DoVyMY/Iccd6h52AhwOHnn8GQ5UR
WtbcAy7IYlBLduisoA7Kfk51QDwzPph0Zc+NHo90APVUcMo/Jf0BMO/gT6imMU7L/Kw/DnqZn0Pg
wIxbS98VpBNeDzrhaq9ZAl7/uydOvqqBkRvCHXxBI/kh3IEgZZKSQgSLs3xc
`protect end_protected
