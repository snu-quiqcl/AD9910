`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
S5Px4cytq8NM+VXCV8l8Vk5GBnqhx6KOOws7iRSSiUtO4iwV2qssTWNyVywBS3kVroljIe6Kyo17
Gwyf8IVqJg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lkRLsZb2gpkqSCsWeTB9blejXfDb/bwR1wSnp4udGk7lgg5yonkPqtNk+Au++fH3vVBpdEVKxRfb
y0SU8eoSyIyMDYaUipv4WFoW+UKpzGoMtM2Hw8c15B/fL+8lNA1lt7wEPekaCwjMi1kyxk4e+XtX
OUbxCNjIaWCYz+bNE+Q=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MCZvRhQkVdd9nIrwuey7oQvO4SexmaBRu9+V2kfj2SacXYFgQNEqnMlDPEn9DCujJvfAASzXN4y1
Dt5rn/rDQX5JW+SukoPPnQ3TNXQFkdEPBq7Zo0s1XmBLxu5WFPPe+9IhwxRiqbbr6kLJ1xH7NF4X
SoCoOiHoYatdxuYFgbEqayZdzbwQUMqVO9wEK/CgsHrmiEhwAXzp6r7x5KKzcEFG1Cl/4883EayX
s2H7rljCGVZQbLWjOTBBs0FYih/0d2dXqFinOYGpRdhzd3CZOHVVoeJvaUrG7qeJmfOhug9xUhKI
Pumw5iZlq5llHWdC0YclIDp7TCFZefcrbBwSuQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kOOuvuAQA+ijtPmO+o3HWYVi1F8R62orBWbJibjZhYhj5Ca82uv+NiF6nOB8LnSd0Eii10ANo28x
at5YsbqtZh7qSygwsmIg7KlimIvfm26Ph0km4fnoDmHIgny/gpOaqKIGVuTwHBnei5jf75yxNd1/
jzfSWrXh/Bv4jS2Z1mrH/rmvDcCh5w59FzBhtHzChGIXP8+BIa0vrm3L+05See7Wcq1Ab/oqzUdy
Thl30hgvyr1mZj3uarW5r00y5gK8+I1yvak6xmixKeOBKvntSsu8G0J8JgzhOCqaTFd8qJlypITa
BqdsrqpVWZYShYqPWLN4r5Ia84xUTE44Z+G4lA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EcdkPmPIpqjnm6VEo38lAHvTXTCOjaJnnXpPc8z5UbFTebo1QEu7VLAyfeZ7NcYMGg3BYiF5hXNJ
DnZaCmxB0TMQlzBfU1r2e1AnAJxMFdY9t8+tZFKvCnM/TL03Y+mPA49b9y+63oofB4K/mopra7Wz
QYaPTj+HRenBQrLztW79vslz1weYN2rZ3+9zN8meOiulF14Ufr9cEnF83RymCa7+6o3uTZhBHb98
5rJiwC+zizYVz287gY/HDLLZjfGwmCCS2qibTVfYP4vV7yWkeCprkdWT6/ki0DrXMRmFMwpZ81PX
HcAMRQ4G+SXbMh9tMxmF/jYOs2dmSmU84JFPDA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DN2rhDPLxDg5WK7mLruyYd5tiB0ZUf8X4O3+oxr9OyJ2QwohmRlJODBLZjEpOS9kzCDWfFhPptoo
3m3aXBH9DyDrI69cG7ySsXprGiE+Vq26iempd9BY0q8rBUbUZygIXGeHjyVwyfuymZOM1mxgpV5x
lB0VxqjzJBYqBICz8cE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K1RoN8LXCtw4zolaAzMqs81xbL7bOkko4JFzYDYClU7ob3sGw7eHwZ3WU6ggAf8V5b3mP36HXnPc
B9sRy9KsQkNWUkLMT+yi0ktzAtq8EYmBKPsw3vFwPueU8GAAvMsMHebrOWBoF6TYabb5PTcZ+2+0
1y/6dT+rZ0PeiZgoB1+VkhxiGjRtWcL6Z6wwR9T+R94pjezzTUHMqMDEjSLJNhNU5M/ztoxgGiCE
DPrSPbai5qfcgykNaNBL/jS6AiNkijwiBbvZ/DWRj/9CvXxWqdtlzJ+PNJUkvl2bsildSuyEnPaN
hjiMhLzO7199PfEVWgqBtwDKyhvOLMjlsdpyUA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
arL4Dyl18SkkFxm52RPRfUpxIaSAMbm56Yigaj+J6z1Gp/HtrgAWMsY6m20QFzLvdGDbrpzbVPns
qx/yB0muMdESCB4StbXzvy36qKW69S4l0h8+bUbFrEAh1hwFJe+L7afQawi6PMivr71XhD3QiDek
QQMefkzgkOKQvp8+AW9AUABmHRGQbpBHvIZ63O7hJu6uwdO+5ynrFqMwBXk5TSEXt157EunrGmIH
SN5yPeCyp/bfxa/HL777VoEob05htAn5PVKI0VtPcoto+TB/PYxppoqwLwRCgiyUPpDZXPiGsil3
p1jqifUe2m6UewPbeNK4OnzcSNV5fr4OUIC0QZ998YZJiRv5fIZ3eGL3PtTnQudNcA4hgyPzx+PK
u7BY5UTFpHwtPtDrRX36Z75tCS3+iFplNb1s9yJoNkRQ5Ut/vStX6smUP4b+Judd0DLcWsgT49iV
vumI4KX6EYwwz+3KjWk8QuDJh5/r5LkmK3I0Sjmn5PHs5gI2hI5ZaQk6eDSp42QwiDIwQ0pReaUM
TYWugOwFKTxJ+FAuzaURh4Yf2NoSIyvNYDASTgt3X0N0PPQ6HqqOE+AyQTc0iOylVz8ajPz9rzPL
h4yt2+nKh4Fa5557dQ90jPSi1Cb+wp/L+88bUIM5LfOeSguYNTgqGBIRTgWHlAAA5l5qiHDM7+F1
qwsUGdPG0MEJuuPwx9PCgHvyh51q+HAUM2226wHH2o5Nog8TuxTq9C6KIy5JsFgSZNmhVq1tiiyT
33uHrpEtKK6PD+kCHJKxOn/ukO338WFCjc0kdqLEGAiD+Fx0Npt5N3BoPmTQl+pS3Iks1bXe7sle
a7PAeEUrgd1wvs82/Vi1ydkjJc8oqQLci5/K69WuazsgT1qxufyn6HXk3uxEDnWRbPcaGABsUp69
QFAtQ2SnP21rdY6ED/avOAwRt4ircma5Pu4QT2eNaF8jC134/Y6y/D8yExjj3QvZsVp8Ga2fTzJx
F92MqoWFjCTMDXne16Ddytrt0k/ILdDpXnpHL8P/ZW1/MnrUmE/x2G3faPe+M2/AjR+ZtlLYfkck
wN6Ry0j6FkuuK5tWRqjIa6yr+/SZxNQFlNk8nMTSLWRiXIgDtyZULbmz42sr2ToKfFVgJTSowrrN
rGepcwF9JAfRpRFPCK+VChikOjLEEzKW3ryN8KBIMkPUs18HTqoMQJhLCjIeO8RWcEbRwdcYRBha
uYzURUiWGS9sX7+C/wn/49nXx25idqchkeNPLmx2b6iMJ47hH6ABsIreE4GYXt547RtZbweZ6qmY
yI7JnAYzuBibIGLMyM8G/rrvgsa29rHl0dNoMwFpwoS88xohSl9Bv35ho79IfR/gRvPpYfN8e8hw
pGfp0ohTgXEii27Qa50DKsQpBV++yZp2s6nTd94a+FwPeqwbC8RxtHdeYqVJ1I7VEGwaloXsuKNe
GsBPH0tB4PVTQ0sXQF4BvWFr/5eKrbbZAbzvJpfy+mdUiO3s23XY+V5z7ePAVEG7yBEY5NWhB5Cn
JxUqCON7AOVgbErhotTkHdlbvNUgUpfG+7rGftBwgWhLsICUIpKcZxatzbeggMCSpvsh3wa2shnG
fIx887L9jYuIYcBPm88wBTYp/KwPKoa0ImGVcqbTCrWeXNsjbuvLHQJt6pqHrDL956omR5+3rp59
xqqQ+2GkyoA2a6Mmk7MHKjfLMPjNcjnpN9iUfZNREgoxn4kuQMNzJWG00eBKhHQsfIX/Jgz+lztQ
SFrj8gvgZCQnrDHwnNLQlEx5DLxfCH1qQ/t4OUoA2LGs8vl0YCXFF3EAdv09muZCP19+B1vTJqZu
SDhKMa0XINnPdFY5WWGarabzAyl6rIL36kpoYbjRaeasDWlSsFSksBcJ/mRRZnI9I5Eci1T/mWkP
b0mMMyZgtk2Po/ripaDt1VFBTO3HrgU2i+gsd7a+zLu08tASyjhRpNlqGJ5+KPUFDjUMrRY4RQLu
3F3C8qdvADfS2qWDlTFr5QuYym7DjdMotS1NRTBbkZUm6BqW37zHpHkJ0gC2DXhY/U0uo9hGXWlt
RpfkxpEXrXdnet8uICekXjHYPBTAno6sh630RzdM3hdQduikJv1azTrAHw0mA1rv9SVLIMfxB6w7
vAcpNEiAWlex6BWwl8TKhQUaFBXwWDPt55PMuQIFOtygi8SjiA/CyQ5WQqZ2DICyf2xqsnVHYR+F
nx3S0TMqYif/Mqqrn04GeQlaksfO5j3+3zg6ZL5L+jpR11D8OvAtuO2FHHdTfcjMpzUfY3ETpQJM
8HdgbblIDciQ0WdIXQDVAw5qZPenztNZXgAot3iW6oWU+m4hyfasdwhaQ0c3biSvK4dHqzF2EaDk
uW0bLqKH1o3OtsQ2w/9kwWrPTg/PFl3Z8vCbr8/GAeOEijpaP8WUhhdVVlcIbap9TUe71AMNDoKm
PyeTGnDeg3DoCxg9kyjUWeWO0Pvxrik8drwDJaFFTeD00McON2uXACpCu3yyEbkadmwElFO9JNnz
XOl0AeBXw5Vk5E4lz6A/l0ZHe4dcz2Qj7D1v/RzyOyumI17W9V4pSu58Fc+NV3z9M0LKiZyc1zNK
dEDC5PR+WuC2ibxg2Mmlv4G8t6sxSQqRgh2mtS5GEuUAN44cHYrGzeksbV5oIXQOHunVDIfgAlrY
qF6uCelMI9han5AvA3WG2e22C+20xcohGhUr1BTabU3Na0p17bSTEkxLcsLg9Ycn02m/YC9qOQwS
xKwcA+pbekl2165tEWOYJB+DjNoV+JPb9BZejtcOwP8KIHEGodyWVdF1aQj1FP6adti8K+zfAbHD
X3STxVuvbqLLOkUPZBFBRTZaiBV8oHS7u0w52BWlW2KqMgEI24zk0dqxePtwj9Qw3NqJjRgbRN2H
C5Z/V49PlshtunD540eFyJFWqy+VVLWU5svyKm00K/HEllByf8PdOV4DO2ceSb1xJUjIFaaO4PbH
rV17pNwstqMWMOhmsoZTpFJeNMVP4+GHZamdmRq4GF/97HYxg7UCRO7EKZk16S3sBahF6gUmp/Iz
34zyjhKJoIIs8pu3OPnU5nKPRLjGdFRnZWjTf6eY+cyu+a+NGHQ1uEKxsP7Em2wAID9W7HI+qeg6
2Xzqyu1KYglXLOEkCb5H4dQpTqTtf2Jh4bfiOVhQxTP0XU1li22wWfUi8tUPm+Jf9EN0mkLvHMsX
eqXyvXAuDuyg3XXxPEi8Nrx9SxM3cDSsnLwbjAnIvdlhiLbzykFUYUAlhxN9iSaP6oForEgsT57e
ImhEHiyjFZZmw4ofGHZqds1InMd56PzmCQHZbAqjK3l/FaoNXqTiFYY/yl4NLu5NAzMDC6vJVB3y
JlS9ts2foP1L1vOoVX6Lfcho5phX37q31IeFlgHruwB95SvSzKqGxrx0wjum1AE1JRnXML1NyuRe
Dp4G5E9Q/xKsyqmG2JBl4I8WJiBXwr81Uk1hOHkEpQdQKVS6vmteRxdZXvaUyqsUgKGJGK6gk7fT
InwbYWwTYlVTaz6Y8ID0EVCVM+Db1BTfhbDbbw47ES0Arzu/0NTItI9PXoSF61a6rVt4rfEpSkzm
y6ityaGpZOkkzIxtrctlYcZCtl8J+i+ZWBgBB5rFNur0nlv/ORkImaXmL5cgGfD7cI6X9SUtcsKy
HeLvMoTytn2jDAWP8Nhml70RrkFxkOfKyFKfCZvP3sQeYRdMSY6Yf/5yhTwzNg4pZjVgXVOusvGf
1Q8kxQTA/4v9ythS4rExODKSYFvHBMAIeShF8CFt5Xx5LYhE9ZtGNNS1LcQaRtx6Lxf3D2cIL5Ay
EjAY6bNx/ujZGmeUJvzvmQW/5EaR/pdqXBoUe4xYTjodKIdyVPbHQIWDJtyG2OfaV1W3AXrLDUNx
1V2GrP4XDRJ8AC1r8wWvIf4Ubu4QqLtUrPCs0VuElL609hTqAEz9DLQ6zucAjAxIvjPK2TE1pGmL
7FAXs+nX2y5KTKZD8zPV0M/nIwuwjtqpkXb3oPaQD446FOyv+q9j2odcdSH70KhrX4/z0MPPByb3
XYaZk1EIBPj2bWdsHtp1SXz3RcLbog+YBtWqfcIFLZssu++zm5iVRycJ39jur8gp4qIRT1Vxt83T
8ro2RWnfMpEelU25utNNga92dSqMMGUAGLZ7M72sva5uxqaDlErOstUekL1d41EUrcLSjJisNfmZ
WNBQB6+UC8EqtvMUhLCjTkzIfhTcVmkVehqXt7nBgw0nO9+5cUCHSZcWJN3YaPywnx06KXgOw/Dh
IRP5/8h0mnmPjg3MTerJ4aR+b10Bsy4FqnVrx5V3Y61Wn7N64G3ZzgVxwQAZB6kfa/t7JpY4BCtb
c3KHGltDO5bC5fvYrIYgyLUtm8moBM4AQHRjnTw40Qstuq34arflpi24iCYyzmjv1KXGMhwSMkyM
VMyN+tLL419fYxkY6g0jsVzxOEZsoeXbiUqWWqkwYYd1YsWleDxJ+I5Q3Wk9v5rICh0SRprwWeXG
G3JHcQnvAAgkb7mdscQ7bmlqehQGLbAQOuW4cBvF9Wag5+QVWcKI+rIwuaR9bRBcLD/D+VbVfu++
Jx2d8dtW4McXp5lGIacftcBRq//PeqPEAnHuMq0l9CXnnJkzvoSufVdGDEGBC10gVSKgxzybWj2K
AcpCe0GmViJXOx0d+KE2FokFBYgVZ6Dyym6Hk3BafPPXLGuoQsmQ/YNbIsm0F+YtgJlX1SD4BV55
4aT3ToQspFR5XB4tA/WnP9d4Q5IdhXou0WeCJA7Pt70yOS79zbBOCxCUvE82WQ8Muv71P1KYDDx9
0RXaN8twBeLiEpMMlAp5Ik6GybYBTk+xRfC8wb26He+Mvu/EUTM3qVF7FT4Z81nKbi8lmWF33/jn
tApUv+YYgur16hhKghc88T8Mg1U7jcHckykYvhYwV4sqjqHygO2ZSYlaCO0i6AvbRc+Nl4nX3b6X
CXXoA5lbV7wPocM+00BwWIp9ZlKzB5z6ldQWxiM+1ACgR8dMSLQ3+/DzX8sxb0CNm4DrEELHMU/e
PfJmppTX/8q6tBiCm9TIBCFOCXUbWHGJQ3eK29Bl3IffaHfdjRwF2lqeWWbuuG7YvGBcshgoEEiD
kUnGQ2MdflYzfJFhyzXjhJsQ00Bb2o0F7ASmH4k2nA1V3m4V3fVv8mg/OmcwZsnKIWaBouHioKIX
TNm5/S1QAWG9gTOlLOdt12Bm8jsZt+PKsBxl/d55B3rZdyAE4+mtqICixUfJXJDs/CmjBMYdYrrJ
PuN5iSW3Ln9X5ZDTPl8t1uA/JvxstDP+XZO2Zvw/I8BAuJBmLGpP1XAxhksDf75Ow969e1VAxhx/
tGogDK/iru2yBVrqz2L3EXTq6as9tpzX4bvcaVvpxNPv0mFQmZKzrwTA91pAdTzrjgZppTDNk6YR
EmWuskd+212KFPti7MzX6MWwMQNnVw1NXtwiVtlK7nR5EBiYYMqdcI4zU45x7nZESUXBWXkJT039
ik9/zRq6uqb2f+bg2CZvzYAL0TAsSggdNIME1YpNfLxhc2rx4tH4vP8Mn6cCPds+kKWs4Bh29FMc
ZpZY0LM7ffdO90IwmK1VvMHytMyjCkgSfiHDU7N3wfbqI/CNCMSWLX/QfYhYKo4BdQoX/EJzlaRQ
azPMWJqMkNKp9VYDYXT/KQdbmumqfPCjQyReX003B8H0cbotex9ftyfvxr8NhzuguWRTYyljOAqu
SMo4/8Vselgr1sbCCHKP8NPCGJQevHwYokX0uWcr2VQOXJD9poJGWR4QccxVTf5Cl2m5vWyqoGvz
xNdZgLddD6cV6BPo6WVqnJKwa8vEuSCvie7sbZQGjKbg1brn36zfzil/wqhgvIidC1fxmdyvD78/
OUd8v02AFKZTBac5j1VXCGBeumCtlA3RKtlxDvTIq3TMeiVcSIhSil40zQGg37Q7qiu711RIqqnM
wIKQMdWBz8BScNeg8zGSt2zw4AVmvhWlBUJUi4VD6gmdWpjRHqJDo3mJqjD0Ocm+qCFVeLkcRST4
sUvfxT4/047IOyp3exd/dDGqwXtSM31JXC1CNKVMVwj5OYGtV0mqZ5buEy1pZNrZSpwMtaSAcmC4
ZsuK+JDPzm88a7nu36K5shhJAgBTncxDk+qx8jvYc8uNRunHdXQAqm5f4CMpyJpt2J5sFmTTs2mm
Oz+KnWyKIW0GJeM1jB6F1Adk3CjK/y5riMpihWAw1jRYEPX3LgLR7LbFzaBdw0TCtq1bbcobU3p1
b7WbpUr8vqW22T06SP4BoqGMUk0XCaDWP5mGI4L8/dBNuCMOth93BChwpugBvAA+xpaQG/RmY8RD
nHwLF1b1d7q8VAR+2mB86wjU3PX7XRajWEgZ3jX90qE/k+pR4W0Esn4mFD+lA4bqCzxslV0vlJbm
O32I7UWuC11Cysb4+WPejRG7AAE5ISwO7BtG7to1meRwOSQ4xLJOzcLHG0Ypy1J5GxDpqglPRezP
T44t8lVWH03GNkIuipNe+p15LqItgGPJFT1hcr6qmM2Ok3hnoeiVOi44DxX8v4FriaiLM0uAoij0
399yuvQiNlGtrVgqdGZoCf77dbEUFvJD2g5tK5c3t47AVasUDsXGwWOBR2l2OjfEIyq7D3zKWS31
dK4enwA4Jy+PrHh41wKm5et/Q6dlA+sSmLzR4OKNTihKT7i+X/BrKUzww67TCfBZ2wb/Tk6KEB7X
VzpxCbwL80MEzAAZWH4o17wTSqYxzRcY8exq/bvqURh2jX/cYrCrJwMSN9gfPHjOr573KGV5wQPT
27IVBSupjfkIIf/W+xLMVajXW5ZkTJyoZZD33fJb9PimP5ESuLStfjZPgvaAGE9UPX1ZUMXodtMW
H3Gve38I+7VY03XuNx6LdNZ79DqQWL1wG6XH08sR63BuK2QYQmpUmsrboEiyj7jj3jOyOLQCdmB6
EUbrFpztayQ/+3/UKFV/rbVs14q1QlYUqXC9a3COf1eCvwPWFIQxWPaxPzWna7yB7UIR/os1qI5p
30CUckJfvT/4ILLeQmvt2pmiJhINyFQ0CT2RLx7qMHbnMhFEEq0nTYrKe8FBD5urSTB/4IuTT76S
gcxj4YDvNjQhTUokxpvX2HlbEaEcGdDuHKBhwK7Kn2WiZ8kFOZWDNcDiZX0VoxC5BtGClFQrsS/0
jtrydc5sIBxvHHi9H7W7jiDZ23BBYsJERGon8RU3i1C+y6avUj3EQgOd9tYfRo04Uv5JItPcqxDP
WhpLhZODp81/yzuDCEopIRJ8EyEHs9bSpSPfXtH6qTiIDpCV9DVmvB+PORawT52e3lx0v89rEQ95
n7iky9DgJ/Mtzy2lsA4tvINgODtRwRWHcigAj+SloYqX3WpO6dnnM7ZqRYSDHEKkuGJbnlSzV9H1
0GNEI7EBD3Zv9dtRaP00GW8XNrf8Px2rgXLTIbsqElasnQOawKic2UikJLZsAU1BYd62iLr/lS7S
ZMC6tu2bvb4FaqeZxjIYYP/0welkjeGV6GKKYC3vWlYejIsccsgY+hJFTjWFvs0xwzEnmTBtvDtj
cSAaskJzDOTvuBRrfMLnOb2jxruQ6v24cZfafkqigMOS3bh2zbfzNAOi9Cy7YiSPvIH1A5GHl9fp
pOUDqjW1qP0Zq3jNDbzls9Nwl3J9iFe99OS1aQvjCyuUB0FLUm8T0QPjp3+gm7O8/Pk7cpeHBVcl
LMDGfs+Rv69SzWmo/BiA4BSADflR/Zc1gsRriD9YMIBSUVcR+we3HpzUDefDJphyYsd3uS6uGYKp
6elz9hwlB83gExku4OWnYfph7pD9pAajgDMJulp8204d327ugbLNp5ME4FmW7yRFPsISj6d+HXXg
i8P62avqbQ7F3E/mMG8A8t/B+oP0dtwYzQoeC/qZqk9rVeuZkGb67qsgkI0TxXXqhR49l0r+BNi4
5tSi3geav3L9RGwVIv5/Z4BxtAt5Xvg4BZj5PawiZDq4MFkjY4AQ0BCQbxm447lxyM8KKgrqZs/p
+arIgH/l2lqCaVPvUgjnJxZo7JCz7p08ToK0k/ZxoABpLgcGVGSysW4yfQYZYL2xn0DHbeO6AneW
m+zm9H1N/wOGN0FQyk0pPED09AcDmpKI4wmmpK4lz/PfkT2m0kTk3LVs815KgMPB5Px9pqwu4ZYm
rZxohsMANkfuXUmwz4SjlW/lzzUZUENmy3WwaUEnnmI4fxPZI7FTqO+XaI+53trN5IdBSemXgBGp
4D0116mC+e5S0FuVSasGn/NnlUYfI3UA+V070+yaPQI3L93PZWB4Ba2XRTm/atKiKkHIivpIQWXJ
mWZCafDxTpWUCDzwrM/ANm/aRh4g5a2RkXJ98ymuK1id8CV/1ZkgNxXNljQ2e6Ux86HQOPdZQURZ
IIc0SVl6TE+Jg5C5euJvXUqFU1m5QXzh8/DPFhGcy6XCoRIHEFDYKqGRmD04+eBFT1e6g9pSzb8Z
xmOAAejsoRcq/F96WfUWYK11ttAcUricaN9lWG5atomhWPzD1uIlnzQrtdLFsRgOIa8HU1rDEdC2
coNzz9AgaEUD25hAfg6zsDtXJAygzS8uKX2/aZVI0NFH+CQf7Xjwo9SgTaiCCWNVx2imkvNyYNpI
iZ0Ysdj7ZUUBpwRXHiZKL0DdN1BUTxjSRfEXu27NV5PlEYopCJhGlyFgMI4E2ugIm2PGhVU0ornT
ZTcJj3dgAE9nan2TpEEoQ6fSLdFaSDnSAn9tc39GCMTbSJCtEVNBc/9wXtJPCik/n28lGZwrkO5w
gawQBeSj/UwJBgFI5ewwUv+Px7nxX25lP4Z9Vh51dRxNJAA4QtGmj/gAhWFmIeh7cn1t6g166mgL
WWXX3HG4yNqUel/sDKOSU3WPjtqUadiQlG+i+/gLYiCfFs5NhwC7IaeNKLoo/iPNh2pZMlTHWZk4
yRPF0CLQAXeQSpNKnCGOU7F0MG0pTYBPHWUVtGQ8ZW2vhiFcynBmLWN1IKXLQAz0l1X8uFbN4Ovg
w2shAgdfj5/rN1BNDqbI3peOLZUaJIUAahizd3bz51JYQ3rPDfcKMINj3AodfQuYSErrAFntoeve
8I5ew5+GKGav7EXv7FCRgewPSdhxorxxBV7rlkyJH/3DeRGqDlZZ5QdkMZ29PriYsioIxiZPcPUN
wuWCEdCbqZxqw5aIbr/mUbSKsvNtgXVtr55DbspVIYPjz2jooZw5Kzb5qQAHB2JnBQcjJVx0bhzA
WI/xlOM4efW1wGxI8CyRYBJZxtnheZNWZ0mBpkGK5BsEFV4Gnriw94CMcXizMlGN4WwsExNPS/ZU
mvVIN//m74viS4XgBwpFiLpblD6WsLmEloCnHQvl+sdewVOZmGW0XmrIaDNk22eR3QEQmGhrwN++
+xnu1gzFZdwk4d13UNcz2PRdgNMf57B4hSffWyqHj1Q9tAl/6D3Y2iwH2LXQTn8/GIGrcG3VTEH3
upfBUVs/nsiRIb0kQXr139W8H9JF9FTMisRHbXpdEZK+FfiUjOH3Ym3sbvQqCwQ8iDCD5p1zw+mt
v7zIltsLZ2edVrp01l80uPjGRx6nUZOdM5vTTQee/twjDm/rjbRZrRKGJQmBQs9xe9IN8rai4s3t
GU56ejSzIMVr0OmEMObX4h/PV062X1hSYKEV5AAo1e0hS4j5oVaMl+ihVCbXxFKZFsbSmbCu9wei
0mHoizeoD4e08NKYP4zh+Sw4if2XkPHJerznY1QJNcdq9IFugjKPf3yijl23SXeGGLrFiaWaf3Lf
u1GxJwOG/BZuGbgYeua2XWvVkGVbh3LhZMrCVZvvHFgwfIGTb9Sz1/DDVcY2oTr8R/AR8QniulAV
uRDd+Ykn/IVLG5CPGEF7ajBPB1LF6HVGS1DurF0TUn30xkyPTP2Zi2lcFFHy8ypEnv7Zb1qh7O5k
FTNbTwaL+LGBpfE8do6QSkvUNU5O3GjZG7ZrqQeaVBXntn7iVC5gxf3d1W//7ZnRKxQtS8nRR0Mg
A0l8uowWCMOCTwdzXx0/7G7O604b0TOrhK82uCH1Afbr/4UBCI2VrINpl7q0xOn1f9EggX4MnpN6
NzMHAW0WLpPw3pNTwqRbgnWiA7G1Q00iNfgblGn1dy8TWE5PKGRYnVEqbzQm4LurojXf98FqVHao
mZ8NnkWJV3Ed3u90zKSEyMDqFw8RFuZoqzJy5+1Dn/NZ8KNSuMv4LnXCIeuHIARENpHUVdtIN4CN
FohNMizyBiCytw/d4pvjSGyhobphhwejrw0H9TxtgNSKwl9M5dhp6kcaOvpuYT5aW/owUcH+htZG
7EB3I0ah/mjOEj60g6+7synBojtppmo8GpK4vIIh1vYjrkI5XQgLFbMpIfxzjIcoS48LVsFCpwix
1QLO8HgGGzesUyFpNZU/zHGF7ZgM3HdZtpBbh0NhvH3PeOMQ04u8PEtCfOsgRM4Bw+dQ2s1jRxGd
V4ehZJzEVY2dfhFnFp1hlm6+9ZbEIvc7rBu5eRS8QY1Fwk9JHgb8DufSui1Wfss1AEICSVkFVv+9
PUx5yp0hWHCjDcTtsJe5OYiBMaP4zO5MY5SfXle6V6JTHwEGRdl/GLv/DRtwf3c+fNu6bJCRVRMO
Dd2GCYI/fN6Ts+CnCD5fe1m8RKvRCof/jpA0VRAjt4J+mG6MsmnHTaxnhJDWm5E45KL+nw3qhvf7
K7HsMRw22FgHYts6VE+7oPNIOLnmGg/5edF2Sy3ex3572VRe8KJ9XwCGcQbrva0Rr638z3QmREXw
6tnw8WkGL2GFXG5LYExShUBL8uRAeGD/svUo6yPqYwZ3RdL8sdITAgfZq8qlD6VhjR6/S9XrUvGB
bcP3Pby0uvUZykpb3vcVAKxjz9eYmeFwU7/SN1bPV0dkq9hQ4wk7gzSQSgB7oPiPrE8OAXaaUMq8
8unbiiMj+7xvZxFpQEhkaUIwIjMFiCqmg56ZYigZtUoqDDtRIluCcKhxWZXYL5TxfbFKZfpMOjEn
ZeF9fpUQz+G6RmIoLJGW/y+SE8reOrX5cLVlTFrS07xlgcPZaimcM5bo6dA1BlsvXM4aUcr85M4D
jCuTNsl2qgJ8JVlrzqRdecSOzUMP9tItbdwVTPkM1xhX7cF5PSeqJuoyu/wcOsw3xtzK3CMRtGoy
xjGJ0jqx1oU2CWLbEicLgj9jo56XGA8gEh8lYvNBnhnk8oc2KTpsN5iweJtMs5WEiP+ZhDa0VL7p
IzmlN5fAhOCXjjCvCRBgV+8C9pOkWgpcfu0fXKC34Fsv38IePXsVreUeELcZ0tu6eGO3Kl5r/jog
05YENoH6o5OKrSFVmY401JAv3pUWZLBJpIDl9pyoMarAgkBQQ9LTQlw3be+UPxQAYLxO//pWdQaT
et/W4q1ZLW5oiSXWUh5Twq+M+ykjpAIA7CrwCc+dsynGzHDhnvoaQtA3SyC+84DaJY25ByP3Ru7/
6+IROIOBJDCeWysSdDaRwFvQy99dZNfcRYgLf2+Ro8g+E/ZSlUTFUYWkuBv/VA+1nOFKnUu9lN8m
UfRZ2qqLvIQv+nNhr1Cvg1l0SZoleWB5OKcj7rAJ0mO/knJwKsZb/XKImx4LyR/9ciz7MJMLQWpM
QIYP9otRQY1fYNY4m6LasrNXY2fw3CeeUjxHKA67ki3HEOpBmsHbiz1TITnukSIkOC+mfpdDdYBD
o8xEuEIZulySf0gceTMsujKXFHuTGUuxoulDYIlES6f9yl7yTeRmmuebeY3oM1PBkRJ5low3egkm
mt4ZbayHnWR+kCvxRktga71eg8qzinKfEfsxdYKGA7OMYwgf0Gizt5fSjSv7ALavD2cS5m6J8Uo2
YsNGPpmm5YGVAFu9VBVwZLEeyeKxtPNtCu6b2EpCH1bzxJgTASoXnHwzyrJ1rbl/LdBd7yDt62f6
oNDOVM88VEu1FOXfeKE3QHBklDRWvtdiW+AQXwdduxqq2ZF3VP5Y4ll/+Jd8rPqz86N6xlxlSlnN
FfbHOKaHyBlIs8IxHwTuyMqevTPn5VUCSeiY+dHjuKtFzjSjd78tOsj5nICgQ37SyxqLLmbmUdnA
0gAL+nGWUnaZ1fkYRVN09odD5UMQroZd2Wh2RoVcjbn+FbTEgeblfRDgiTgFljgPxxiUbhuUdyn6
LhxI7JqAX4MPtzVmfNF01AxRoPFycwToNoWA8cAbugXCbPoJjp55F1/WWa5h0j4rADZJZT2P+SKd
eRTJS3IH4jH8+Oxs24TE56Ygbe4FrxgLmEutoYuVHFiunUa514He8yp5iMtqcNyit6AkhQqfk9B/
dwYYn6oow7g2LlTccM7MQtBZxgW2ZzIv0aUseDqr4JOztdsfQQSXci+ZE3DM8d5D4L/PeBWKNMN2
JUzFCGJ0gcAudPj2lJyCJhh1N6UanKWx0jnH+pNR5aETj+ALO0K3J9J+KhsLMuJkrNNmnoAjYeD1
S1NSkq2RRQuGaL191XptX5Wrq8MwZXsZ4xKPgOOC2OM+MRE/Y5FrKVvM6BQ2dW1jWrc3IwVWP0UY
XtZJTeHPPLZGAk/5iQVKAyhLlpDkwsllO152ZrgWqeRku/1jzes+ztpCvtZ2lx5TdAbu7jMUJqlW
TCh/SAEEj0RF35g6pIithxy0SYxVOg+0K1RR2MZOD8oa+JfuBN2Kr6x5JhRsVs8I3lQRj7ws1oEb
n3hNqr6bw+aJikMBsZAr2ba9YjJ5+gAeyQUd6EYZtQ6qVewjc6FW66odEh38/KJDlMIbSxauXu7W
P/IIYdlHP6Pxs/uMKJq6T2/BCtGfwkvvg6a1kqJQFU2vbmK0Hko11K8tRC5ilP1GRJTleVSMeETe
WJjFVNV0lwgfWDingIrG38JD0PXiIRYgQg+2LbonvdNACKN9f3Qzw5AIY5KA3KO8Pl73lKMEQLYg
k5VN/prVeFUqu4w67/IsWIiJr8ycMeKXSJIWyBfZYTWXxef0CNDCMcBLR/W13x7bvlQhot3UnKGj
pliWaePR1R+Efq9dLWfJ4Twg95N6oGrZt8ufifQrgssKPapN1Nn93sXFOf+Fq//y4ta6WQOg7VWc
9g7Np5CUmBreqe/vFaCuQEXkNmQWUbeKAjXG446dwhbryR3wQSReYKoK9KwXfsh4U17oade3Jou7
+WIbUJyyygazwH3TuazZbZBwZzMN8gyEUgmlj9JbTNlBKL3T/Vxs9YSHhoe/Mmh54PDmdQu5fuhc
8Zvfvx/w1AUhSSKERIL4nw8tTp85T/rUg+s2iSQQav6nR5jO56MzX7wSW7lErgV9eOYKgPGOW/DX
iKlgGcGfOeyVYFYtoibMWqDkoc+6ieRMoZ1rfd1c6jSwiVFvvbUWGifKYnlD80YIDHd1uM3+MDdJ
p9Mhaym4xfgwqkaA9vC+WqKi5R/JOOr9swRtd4+ThyEInm19+nmMNyPUsp6+WN7PZ6MKP74dL3vC
5noeSAz+O2jVlJKBde1jUr03qaIsf/9wMSqG8ugvAdss3wPGP63yL7MkMCKoPB6GgedSy2XuHX2d
HyfmmN9GEcPKgKAF8KeFWant8d2rDLLfq0Ut5x4uHJ+Pk+Kvi9iTt0bNVZp4/v+pbfsKvFHI9vM4
DRVaYgxpBgfRrYcFjHOwuhBxs6rOU3NkcAR7RMHZ14dTI0iRxc4BSxgRWP/2q8aknwdL6FC5umL2
VnmsMX+Nnh8Hkw8Fypsy1mc0Xl1BfdAoixx86tiD1YFvoYNYZKRJIujodDUuxABC90unKrKrlorI
CWMGt2U/UHPnYFkiKPfh/g9HR/Kn6h91JuM5hlKEVZmwKKN3O9LItNG6dhFjTkJEmI6ol/GSMN2W
853VleB4vxQ0cs0WSOr4HAyqaQBzXkh+DyvikCmWjjiLLZUzEqbzPX7mZidMFi2hwDfRHSMnWFj8
U0lcjdzOQ1NMDDpQn42wrohQdd5+s/RAJAbWUhU+uclqAoIB4y5R8gIo9UR6/5qGVU4mDl7aVhw5
oGVUQDD9dJL7shoX0Pid8i3OotCsh5j77G6ZkrEU+0jpQBM9zvEo7GGEIxihF/mLw245UM29J6eG
HbG6cN33v4ftyzgsGgyk3arDCqCHehAQ/5BIciGhpksiq88AHM5pnwjMpcToOaAt3s6gwZWLMYpX
Kn5X76PTCa9ozay8BNLec+oMqmfw+L/H1wDf5N59n2SUimQexB0bS2VwfyazcxQ7rCEpui11Fxot
tXpB3/xjO59h7ZhXw83ssY5yKmmozPj/jaqfHkSHA8tI5JqtfMh7hpp3P9AzHD7jVxElx8QkWtsJ
LNKHfFF5wVGPRp59LMavt/ulGOIaG5q66akGis3QGaBvtYzC6NPK0VrkLeFcBp5lXZ1FJr88/yIC
xArKDkYZ1ewdHfxww3yFUz6M4QZfJ7+cAHlk2hgHPnQ3mkrEgmHeF6uIcROK8U8CbacqoPw7FicR
72ZPfxa4DfJ2px5apoda6S+F68ovd9GbBEY0WVJgpfLxtLzW5Mr6ndZeO0wg5meOZ7XPHpPAqvgQ
1GTN0qzPnIkvz2QuKONFu/FnOpwmrWHJH3rR5gWUZaoo/FRfXFmLf9wWbxpG1SLmasHclGqLgkpM
oR/rQtbceH6NcSAlZGsy8cvmDoUTgA616LGeK84/7+Dr6Bi4rmtjw5rqxMc3QURWXg4P5NXyApLF
baJLshc6GwTSSss6AmKRKQBRV8bAut67WG/H4OQCLbKiTvSaUTl/Zqf54vP9hkt/q6JYE/cl/Ym/
Yq3C60hcS5v6hbzjH3gavIm88VyxO/gC0lC6gAyIDOQoo58aPJUyy9qJB1jGtCh9QGm3wGxyxLex
9HyKwoJMxuiqhPuB6IgA88IklvnWZhmQd8las4//IU4iSk0wAxPiRRgXPJIB6p3UMMPIpolW+jYW
KkucGT4NC27kAdaq92m5J5FupluB8g4pSD3wqPUmXkWZdW1GRPLeLyBug5UT/jNebu5vT5NrSjY9
Pgv/ExTxf9Bpriw8u9eObYlKlUmJrJpm6YDfZuUM9a9F3fjhhUqFQYuTGVWVKrGA3gQaulKxBdzk
2g+7Cof4rf242P/OwnQ2QsVois6IqpaO6740mxuC5mnOkEY5G88X1UmS1yaacA2dNtn7eLrQ0cTK
zbiFD6aylA8kgHbhTv0cIQqE4mjCXMFGMIXLUTsU480RSFOXip03a8HmBuMcZ80RZa+6hhQgViu7
zhn4Z6MY48VCcvkvsvpxTx0h6pNa5XA1MLCw45cWEl8R8fzau0K3fgqbsHjtkQHKah8Sg71b6WuY
p+m3hD3temrvTHgyISK/cCCwhwHByDPGKw/5UfkzRQLO2PaJaqWLz6fIMz+XtGyBSnspJ5gM4dhI
GzD7rq7LRzWgGs5V3Al4i/1uqfo0aZg9/MaPViuCIrj9JjE9VAXL9zzmfFsHUc4lJJgT5Odb3MgB
S54doNCLH1IA49779UoQF4YTFW/XTSfnbUBN+IY0hukBzcGCHLa9PCOwqm0LFMt+gmzs/DfFKrk+
YsOv+ACRBXmLNGGOvxBHcyXmNvuDLPDE6vela49mlvs/qS63zhQ4fvan8Ax5lQzZAtmniVLKBYGU
eaKuOJl5H4BdL7WmbZAIJ2eQsvUEDYrT+GaFDLRwtWPmheP2CxKC1HKPzrJjNLcgnKj45HO+mz//
TqZrvEL277NI8X82aOEvvCXXic9cjnnrdCItolErIEqaqMjvIDD+XJ+YiOvqcrLUT9Ubz/LNt9Q0
o7Av0TF3U6LS9QfOS4wHUj/eCb2FTSXZYQCejaG4dCGA3A3hjHmcrEfgY7Nx5bW2csQTVJSHEDVR
ZSpFO67b4foHUoVy3lulQ2CPOQs1QmSegMxHF2cvwcDi/F0DZVOsvaFwFFPjox5nerD/T3LT5XD0
CyfH5zt22Ne6jAblnUKTHfRv5v4FNuW9ui3TvityChQ5BeibA5AaliJ76DmKYtNhCJh8XIreWl6a
JrRoKyNtafKcoAXXxo4e4FdBgAG0edvWgg2c4Z85B9c9Sj94H37Tqv4dF4TFowb8RyZVLa+wDz4r
lZmQUegx3XxZmHcdq6qfs8bMwV/s5eVxQf0OZzNtOenShjAmY/zWgEvzyx0Xg8JaWe+49bZYDEqf
BTmBEc0PdhryX+Vz3WNAXpCXPog26gdJywo9isaxBS7WK+MdElmtjdwilMPNAdE4XMuoE8kaPuNN
hf7k0+yv+B0R3nC1DRb4rJst887Q8iRqt5Zhwsbpbim5dq1NMxOgGYIa/aoRa6HVdS9SzKS6jLQs
Oi84eoLXc446RJVX3v+P/47lrgNlewutp8spKR4QF7Lcf4K96mFKb/078H782BOBhk40A18Oy6WN
7cQhMW0Ag77b/zW78OLuE4VCmDXzrWYeZmW9QVK31UgcYnl7Ef7djoLm56J9GB/J0QIUv+PJhpzi
9tGWdVMMFRGtyrQOYFAAr1zPKCDDryoc1tcNfv3HgfKjQ/c9XJJanuHfV+WSrfexAE070Ob6WTkD
vlSNEThiKAQi6fm+yGpWUFTkh+ygWGWnEld+JhK5Q0iZ5yjQ8UP97pVQ81B6BIAw2PCPC6BgUixC
g1W73NcmFKpwApLK558SnwMuYu6kv6T3j/Jbj2An8btPeUau1m2w+4dNhEkZMH1K2mc9tyH0mywK
XuvUv7rqjuTcekOkm6bkhLwyKJwovT7sSLJEpiPzPyP90htAqJUTg1LRl/GXHU/YoPqrO//VVF8B
SGC8+C41kjlhvatAj/WwkmmiLFsd8f7R1j7gCUMn2ZGuNicC6LL7ZqcLQz9feMAwYY4YfHK1tN2H
xXS4lN7bPPvTJ53MF6fT2H05aTx96U0Rc1M0y3/YGSU0QkZTW7K5t1NnmzyuqP9idrJFzkyTU/Qk
v1fQ+k6CJnyvq7M0p1AnNx4Wmv7kNsIVrMBl9X9HwVW/aQhC/msMf1l+5X7EKx4q9q/mZ+Lmw9WE
OqJWWNYBUPdfu9tGce/wAcDvstCWFBbdEZvlHg0zUX2/4XT0+0LlYdzZWDOFoAP9UEgVLJQObRWG
lzDdJnjHjt8k65QLtbrGRKOzxJaBg8e5+7dfYEEes7TysfkwqzJEUcu75Ei2hmuj6IO/1mq+6+h+
hyvv4ATjEdWZeMg+XxVFwomra4fC6rQaAFyyW6kSjfvCS2YY+GKc4munEvsrJVs0ARuVzLX0sdTz
yTYwaPHk/D/4NJfbq1TxtC8aRgBNkt7EB/XnHYv4TjI2+vzeAbi+2IAY4IwzQeG4/ElwQxD7luk1
UBUdfEXIjx6QT4ENhMPhqfhWNqf9WjL4jt55UksFE0ivMo0hCKbuSJ5issqzV/uc4zneUVJWP5CM
yu/4t4Oswjn3Y+q45TKegwmnAm74xCFuMcufM7cU77QP81ztWX1TOxNrcIlTtP4ydwwJb60Jt+eN
SbXvFXcRVhpeCUQdpg7GvPYCgwGf41NgKRJgK27onAZVBVbBVq49BhlebmHdij0W3e5qVrtj5mtL
0/jrVoY8qDkjainIX46R+dJC3D/HNrN6leU/wXhZJVyuZO3FcIS2Kt10kmRAJjVvY3swE/tCU5Om
7qjwtXWZseqqO9za+qKHUdhx2lllPeyfSreEicuXV1600YYhrhxpU3w0XYU7CHK64hy+tN/nZr35
m/VCPcRKIRwGiu88zdn+6rNA5Xe9ClT88wuIIdorBXKAKiuXitxVejOiiRHQ7iMnbZcNlY7EG85H
Dpu8utYIiPfUQRgaeShHhHpKJW0uObWOTQy/5P1FY4GvR0fT03KQW+EUDP1ZOq7JxAEYjf+ZWyjG
FnL0gt5HJLamoEK/5XahPsegA8+N3EbFdhc7Adsjl7j9kvDXGFIOI1+KUcjzqh7vAsxnst+fsKan
XfeMpYDtaP1ZBhTSpTmY+972tM5ZdKQRp2RCdqmYMALkQB9X+F50QVWkhlV8loYLhOJdclZuBmql
cEpvsFLj5jsQTU7MowGzr/2E74BNngOdjj2jiHYczBngXvg+xLJZf2HOakdwy0PvbiYJQDRYZ4qh
c+oj+pwd6p+QgbUxbOHeTKIfICKfnZEbvfB5agEC+tQxBg7lqez095t7jAMyp+NX8dcisysFJ1hv
AKbT4UcW5Wf5iOWO9tHyodTjhVetphTto6y3GSd7Ej/5YnjVUm+q4uyMV0hfqcm7GgDZBHvBoSEH
TAaLjY5Adp3nodH2ooTaRUthyQyjJL+LDdIYH+m2K8Gbsek8XqBjCwklR9w3k9EF8U5ARuQyYkVJ
by+XlnrCWwGMb3vg3Za7Sk1nnMdRgxPrcvvMybTbqJA1z8TV6dytLQiUPVavLZZ/KnKwPCFh4kFL
22fAIjdLk6oFldBKfk+LnEQVMkSVpBxicEA9rBXN2w4Gy36i/cfy0Z6SQtIW+ogGTLvhEb8xT6Hi
fQHd6ZqYbPK5MbDM1IC0d1yYdAO6vK4pmaSwVEhOa3NjJXNnYUaEnnpK4c3vQLrAJ7ZxroJlRyh5
MgBWlmREFDf1a2yaK/DNrtR4tJ1SisT9ssbQXnBa2nyVmznCeCY9HPFMaJlYg+Jf1f12/ARhmL/l
gpKQEyRQnVCcdkGdb49Bvy4efG1nhMvbuuY0gMbaOBjrR1b1PJB3ZzvS/qLDkodnhDNhl8pdJh3x
gel+v4TQwZOP4Izu/gCDEMGNZHWLi+AeRMT/kuueO/YOI0EcYC81gjxy12KTTFJXWofOcipJ2fXE
H4OCSvI30V/gNNkE9nyVNakJzeBWBaijrt2yFxzBEhi2B9xg7PHQogJx3fIdIMd8oFrEE+MJtruc
OsjC6ovY8qTUCNq/C4wmeLy+c/TH5r4HXEGFTAYbQNtQ8iQujMQ7iSMxr7idZrHL7DP3tsP00TNm
x7YNuh4F2cQVYTPnNjE9RuQwPVBIfVF69XwjS9SlhVlPwojaDB+3Cr6R0glRg7l0v+6uA3SHeykW
EKxRWBnT4PM5px0Sn9Wwofb12B2BJ9gFy0/RPXmRgV7U/g8uUjU4VAx3SWBpGzxxPOx9eBQqZ7b8
DDwnYayaWnV65jBrpvb1fSjTvU6M0Ro4/aIm6N7uC2ttOzm0gEBUMn4f+Bt0OtMnXsCoYtw1P04l
IOLNa0V8c9oHod/riAQoPwWJ+5ABHj89cUaQiPzWD8hZyk2SR9g9tIzHaWZmd20zNUm+PWhfGOSr
6PnbA3fII/33v6r+Exu+6OZPr0oHKycjPZO95I8doF7pVTOfVX07Vtf2ZBxvOA2dLbP13QuEiggB
qgyTK3uoZwHMxLATMuaCrnVHahHdl83wb8k5Y+ZaGtRRc+V6fclVwYmtBbMsUjAlWnBmITpuHUTD
fZVR1+4BPaEuq730J+ZBmnNN5xElTetR0mSQNSf4M+EoFRqkxZVHGv389LENp2oSCckgD7PWZ7Gg
ypY0rH6+ddkwt4nTAgv16GOyOv2DnU6teh9Ygpyu6fg+4Y7qX9WeAT3XP1cNpNNoE5gT5iEuksqq
O9/HjYpoUTcWuVmrZ4d5QdWhrmRDlWZU6MLGbh6N20QT3B4RSu0qd0/DF5hxm0JaCHMw3FpsWQd5
pGy5ZbeRQ0HHXgLEEA9l+dH9c7wdQjWcL6OrdJq1m2F+rHCN+ZZkwwPhW0a98haHXsx6rXXlkG1F
MB7XeN+3ZQd7Y0rNPPUE3n0kesJCI+EvPdsA2unCGZhfloW4RuueFXZ7mEf05+KVb0m+gY+I7b9B
9OYq+LiwN/oJ5QE6bDOr14zop7smM3uez06d3A1HWGEPu1xe8jxlJFq4vphme7msbv9FfuGxQPPY
f4GrrCpqG83UMcFblRad8TtfhsEtvu0NpLrSrvuCZ1zUJqWCIO8dJJIRp3/Gmak2Ns+yqUANCa3C
rYyTBOgAK19B4CND/hzDKZQj8T9Fr1n5EYYk3U0SvCVK8peIpaCCN4r7Jjl95wW+OcpV3+rHxuKM
GfunNAA4ovLdzLrQ34JXdSXNVE2ygkmpYb5IbhuwjJzwYPlqK/bh133PBGP9pfFNwTbOgtLThzJU
4or3J4o7gQGCdwatvdsznMw9eKR2zPrDC611Af/WPgRYCSQcCcTc7G87RDysBaAkF6X0nF1Kszfv
ucJQEWQ3WnotAJTfpCWxgbNB5Wp6dXeXSDLNNXuKT+ROFojFF9sVvhmhbHrs+ofD/ZjMHoAw7LXp
qWZ3hZjS87HRBlLrbzejIrWUA4b235I/GZWz73c8q4C6kTkarxxpeRLoEqo9G24u5wnv4bm4NUdK
CxOZ8tepIwaLa+wgIZNkL49E/EShY2BtxcBxJSRZN3dDpq/ebpScuDRNUPxGQNfCebl/N4nq1CTy
c0bO3zht7D7SA2nCZJo5PoJB7pNN22CmraJhm4FBfknzx3yROyenMrptCq1zXTz902wIF0NnT/ps
m4cFLK2PDCLLEZKQIPjpJZ2+RvJANjp5Tf1vUlluVasNGOW6xR40CDnkmg+3k529gBgmvNqVwed2
IYOXNnxX5dDQOLgLs6sYQCsie0JNJcq02nFSF7YZb3dl+jFXlURAyZBeW/dtBaqqM5KsZh8rXcrh
oIGDrPrIhH8kBOjjLsdQ3OvLoVcnkgCCIIugaV4jtPjaLzyUaV27jMSbo831CltkcU84i1fhyqJJ
kSy9p6L9K1+iswuECaUf1tafPgfcIm9Kg3yvZa5IJeVIt+3Oyt5/tgfghcjFDMoFgQtvswWhoeq7
m0ydO1LxoDLPLDaVSBuOiSCuaw22X/N4f3ZCE/V0yajpq5a+XQD5uuXQR9OJdXwwh8mEX6uC3U4l
iByCg/3tQNgRg8xCbnnwL1lt8Hf3BZB7pUMkFjREpiWAgvc9OuzjYqQaVlBmzKrJlKiX7Ha9D4Rs
VOQ/vVowA2KYNAa4W0svlsRBMFau5+l/1iTnZ41PYmYUjcV5Mm89NNhiQN13MPp6Hra8ZG00N4MG
uX7pPX6xSACfX+OOeOHjTL7vTQ9VSl/UALe1dcdkOzs28dM71S4kDaRWjO1PAM5QAm4Ogl88IrhZ
Va9a4HCPnTsndkKQfdgD70cz7fO1dPqBhhpJU8rppeh/L8hjzehrpKoOg1O0TjaGxzdmpnlYpeqH
f4aIfQmVCJZWw4HKLgN9KzT7wNZaWYolWeEBnkRGXEpC/sC/KdzjjOapL/sA7Ahx2y8XbYMDfNlC
joNRxqEoKEXO0ZW38X/78811KFl+FNTFXcco0AKA76QRIzEUxAsFr3VEyA36IVpBaYmeXlVhMMWy
7uks6JmrBln98GOWerUcGwW9CpOleRLadVHhsXrJisSQArr/kyrbMpkd0AteEp7VZtkTmb5uHR8h
vJRd1PgAxohij2kYXyNKlTrFRI0RMrFLrO1f3pYTA3iNqUoa6c4JQyJ1M2BX8kE4qdLjeKPJFyFx
gHXRmVqVjp4heA6UPCHPdzNkAAob/xK6ruTH3Btn+w0Hvz0UxYnhas4AYYHM+D/m+meruhn9iyKd
VPXr6hoZ4tl3MRqYqURj0jKqG3hYWtVdIFcsz3bwDbNEkAW7Zt86m4/3/3ZPI+Av46+KmvBcc6Rx
MoPIwuGmtdHQsUqXo0LbqXijnZ8opUy6LL8K3OFqpeyfGz3/3sfb2vAxnhmejrVtjPgAT0cWMS3S
ygDg/u1fDiBMBOPZqSkvDlnenRT1AXjikFb58GBsr6ReEgYlB29JX88RjR1oQtEHuN55lL/MxMdQ
PToHGSusim5xw3R6H7nQ6UZtbqPr4KkleuPOZpPPBz3/FqsqkpoW23FxtegR/3zFzrI8RGOZ/oBM
QyvGc21erqskv/9J84QQEW+jEXyL5P8bblDB/xPDUHFP+fdRjRCSdChVDseBvu8XPVHHouasu9HE
OjPMpZK5QYYG2k2cM5fUn8yV+p7yYZv/q13VM7n6jbXK9pBe77N4myMUXikw/MbP4kBOkOHIji9T
JPrD8HHycS8L2PfEPOzSKDWOtslHhdAC/HkeoVKqmXjhnAMNUAwcvn2YmVXvDE+aO5IGM9M7eI2x
EPdn5Gvlqcx+fQWeKZIu82t9pOQn609GZe+Epk/7iF/N0GftarYbybuFsszJ1OV8muDDwyUOIerx
39eFy27GZy/sCqBNRleuDnnJS7g19vyS8xTI9PEfKDZ+AqsINOaI4xtRWITA2o2cW7jZhySoTLj4
uHcX5dag3UHrSRA90ERP4PpazKPhfwUadhMeEQgvG2qB/sf0Opz8e4F4DXA/PEG6pj3Cn8ohRcoI
riA3L/T84MxH1Q3CeZK0oSHgRvmS0+2GKuCp1l61Xa5oF3edndV0IuzBUIY4gMlngZZnbQ0J2WjC
QoNiwwXtgBDtP10okd6p2ogpl7RAsoanYx8YdrMVQebPy1D0JMy/ENfqjwnUjDnCAsoVALkDjheP
1IqlYIco22JUC7G9CWfH7+EFF98jHAZNvNKKoC/j1bSjzNz36VZJnAQwlMU852io4Unz2f7c7ltz
CKR6g9zmiEpzUCOvXg4TaMuFEuphFNdBn5H3/aoAhy5oL/w/cDyfMwHZxVePhidZqtAG0piWfYm6
67pPHsNz4bQ6/0lelbhOzo7M6vqFVmlhmDBjnaopXiTEHHaLzACIxzakRASkc6+yW+jBlnhkAOPu
Px7hsCUcMjtJl3VCH2dGZh/h5gwOAFoY5WZ3B72CP0HWFoLoWOPycZiuTBL8beGaSLX/iXFSBUzO
o7TX/hnf8mZM2So0MxtRE9r7WqMCfet/e7h4lpkVWge/LpfDcbcANlS2VcCrwuYCOwlIEpfO0WOq
6yA/r5xuRYCfaOY3NfwEuakvDErnpfZLrLdiaPJ3oy5V6xKfwRw6dXdOfmC9mY2gM97U0G70/Z2z
6b84p0L7Jdl9KvTIo/yvvJoSx+R4T5+xtym7p0MT25tUM7stTRE7uGN0gOfPAu63279qIYylQj9A
c2w6XwSUAvD7YXByp091Oa0cSF+81GX7AKxQHF1bg3M2yiyylVLVeZoeUS7QJlr6qO4xN/DyJuCx
FGdUXqfU4GzETeJ6v2xXg8kam4BLoMtyABTNvGPGzJkOqI3WBJ58zupulLwSeNkiBcw2hdrHJZJi
a5V0frXHYwBLVlq+tI27YFZHfOxgSZ6KDq1RYMaGXCUJylOOLXdCqrG89N2cCUA7xCUesQyEnJxX
XaY/5aBX4nXZs1ocXVBsyNG950fitD0Ftxr+t9eeoiyGbnbnsIBjgr/9vvVRgBOGtCJ+u407Xwfz
9U6TMbQQ7BSk+//7yuaEFVjwFBry04+M1y8qUYURL18t5AnpICfx1/N+ynQ8OT/3jdF/xnPhtlQ0
kApX3wpK7CAievc+F1a+7E/ge3yi2dr2r5Jg2BBr5Zqs4Km5rvXcJtYGgI7a60VZzFa9XLC1Ehob
rX2pCnw3vALluHNybIzf7gNAmMgig0wxoMY1xPFkEgsHsztLkuVvvkkHw3KeX241eAzTudwxCuCj
g8Hp7H3ozdj7TTDJXDDCNFSrDukJ7K9V4XPWl4s/Qkuqr2ean0C97o04aN/B5jgEfmdHJRVeoYQt
txptakK8IUq17XdODu4MLqXygqW0uGFrGrfGYJeou8kmxgV0W9chbEt/kznvxUkVMX4emPykj/m8
iDbMh6Z6lAVdN4OONRN69koR03WnfB72iLmC+pPj2wUjA0+WRjHbrX6R0XxZZGLG1w1AwLGnQxs7
374RU0HcYlCuEZBHmRTqnQEiOjd8BYWQyoZ3b4/dBvYiAdSvRKTlY1siozBVPl1rwY7+IJu9t0me
bpLQAyDSAvEN1oL4KxnW+TD7KArxnD6VIxCuYAjjgpVuEesvt82B9xVGTkTQ+lfJOCeN3OeZbFfx
9LicyLolR62hWOeNQlhmXcqL23CeNDits+KpNhVhtnjpBaqCrqyP2Mh25qrZkvPeSQIzkTdSZhFd
VsXEl+Gouzugfr13d0KBZn7M2WXG6hyPq/AN0WPcuINY36WOMOujJHBScp0cEFi6AY5rnZnsT19Z
ilM4RcC3WNOflE/tm6jtua8sqZo4adC6tyeHZgS1x92T+NBpaTJ6MP+cEM5WDRTYVi0bazAvwEyY
kuDcixZygrKKAyZda7l3PA7CURKhQFPVZAeOSve7N0xTroP1dRBfv2QN5To6lckekJ2X608eXWYg
3b4dhrAV7o4lyF7dclpJR87Z5NPuvmSULFeQdm3scsQAj9znXh3GXMUzm4i1LS8oPx1GVVX1eRtX
J9vs1xZFGRnwZcoqAYfV+IZLNtPT9KKZAxC9STtF6+5mH0Nh/HaLWSx5GmL+mgGaLibJtxMkEgw4
X/hLClVTb6N239Qgd5UbxJb/JSdBAFRtgw2gUdL5fgbOml/c86b0OtEgISW9lV+lShxwiEalqiEj
4fkjyZLmp3oax7qz2lChuz4k3EofF6WHqNiC274tM9SslIMd7aRvUaf1sQXmu7slkJJldQue1PpT
9YH45hr1eM3thD21OR/hslBIb989tCy7GU1/cRpXfquLddmXB6tyY5VZ6iLJy4ttvIqoaAEOb2dT
cisUZUtgARZ0kaMvKBUv+aGLVc7N/IeIH0kij5eM9i1FA97vdmIbgxuT27oy8ebUf7GoVJ9sTRup
NQRxFKQQyc7/XG/kA7wEBtTqmk3SmDEkYKf0j9E/s0avnIgsamezcKIoAlQbfUNudTAuD9a1lvol
CKQAyi4yCIWmjoopnEIyL11aHGeavHBFUUTmKNlZC1BP74Bkm8HnnyYqb+j8V1rS10A7uT/d0U6e
CPBg0aXXXdNnSjwtUWtURx/qLrURNRyQZOvt+lDcZBijntbW5XKrQoZCkSpCSrFuttztDyzbWMtB
/6HbeLu8OjJM3f0z0gI/Ev7tjPq2KtKycCi/ZCUTh5fUK4IGEG6T5ok9otVXJTQF9YdKqDkmbNJR
OI5qXDkg6ZtNNwYUPyBR7tDzSQc41w5mvzqiZ0De+xD2Bf4YOlo1/0b17UyibKTgfQ/j8bOjqUec
+UqBrRhlYLfJaRfBXSDd0LiLFf7PZTuOjynMaOXfXX6leWNe1zvOplkwL6rGcX6SN3GyRYvk1wXg
kgfd/dLooPRFe7R7os1LFqkXrywELl2cw+rWHlAlFyj73tTROiQNa/AU9/UOStDyh9nD5yA6vS/o
ApcyfQRrgCqbHEhFlPOfI2fz3UbbfkJ6qi76ScY1KZ76znDizG6tplq9+96v+zTGSaEu0SKkc1LX
yEuCy8yy/0YFfHCtoQkh3ujrQgCvIZmn4bwwF5dwfEBVjAZhyDAg5qM1KEqVum/hQJOBLqtcm3BJ
HZ7kiJuN+F5MzpIGKztLCSuSG+pDEdlFrjXBQ5dol3xXuXBzJxh6ybDUVvCQEkNNVvNY2cg7ocda
tK/qG0RnBgYsJEvo4CzjtAJq88z8QbpLEqnad0/KVj0Jq9I0cb+hA/6eptRp+rcdllu6ENpOFApH
NkM4RbxNUyt8V4efivZQcI2vW1yNF0SwYURSciOwT0ghPylKoFolaRi2jN5mLpAp+zxt3sPNgc7y
ObS15iQneTO1eJ+3gfzO12Wv3JJk6mxWy5ZHd4uGTpnOZ+CeaZguhxNMi+5lxlEhrYGxzIrQWowy
qiKej0omMGhL3gKsQU/yQor08KcBYE6T0cahDcuqihrnoq8vjJsytwkv2nvytrGWr1Ey3WbZq/9q
4chSdZKzVck5jMGN8gPnl/npmbpHQyi+i2mPwNayJ89WyAnvJXf4shUhNYMqTzm6CKAtR8KR1q0X
73L135TaB5oPuMuTk3zUDv4ZpIh7QnunISOonD0LT78IuF5cv3G7PP9uSII6vmGtDpIacHu5c5YL
XkXTL8IeVbXQ0rR/PZbUa3b/kbxrPPf0TaDCeEvSmbLVKglGJwhjtWcDON7CZ8/RZQBWhYz222Kp
c9O8f3qSv3UQttLzEi5/u4K8/jXtqM9IFde8chBzKn7xQ4AWxOBW2dua7gXyM2ch56LyqCltNUGE
d87wLWnwulmC1xKhgC/TJ+VQ//67YvtjHjR/+nFTyKoc+gp+I3mnMdfO8M+xkMatd9h1pkitHX4U
QTPLbAUlDUJOuEGS11VHSCT2VIXqil8GA8/xybHfqiYPahLwPyU9x0o41hrN90RmoaNCxye3OHa6
osZHZVpPFjz0Q10vSiEfainbR6Ualtr3O74X+h/aoTdh62B+MSm0dBG9zQ3oVhwHlaIkam1KMVez
iWIpYr1FqRluYnOu7GhmCcGEnsQvk4J2a0uj7Ale1Zn8ChBmoRc+SRV9jR1yC8ZkOt7oodaxPa5K
ws3EvAPmsiWlTtTEQZWCMiX+1nhOBOZxmsuO2qT8UFkQrp29I/RK8O8pTsusIeXYjcouRN0VVjIA
BLlUtxWEG6JN+nzlbDvwzCtbtWtt4tnlL5ukk83aU+lPKkPAJL3zn2T9KDe8jP/TYaX6VbKiVZIT
yQBJPXcG9IMYTW1Ek/wWruw12x/DvVkR1pLkYQfL2Vko4XJxZb8QDFtzk7VeAJ28Q6bnonRagxkJ
2CGsVJkO5BzaYtmG5zZq/HvjByWBkWKh5+TRjjtpKs+9qZlQj4LwJ+M7aqOxsen2Zed+O3VxyNZ/
QSzxhN8A4VdisSJvRFiO5/s+VK1T3Bvx/GD/fFQtGSsLG2Ft2rgSL59yVDJBP8LXxmK96pj9eAib
q1Rt8ukVhOuzk+/w9RbpcSnjkl5x+NV1wC4KRMcF2zYcKk0LGK5/jMT6okXWoJJ0gNm8MWwG8ctw
M6lPl+6VdyqrU1+zmG2CO8SvX3zlSoyhZxYfD0DWsLmwsm2jZ9beWCjPPAjwEWZJ/Un1mNPaahIb
ES5AAZWkGlk1bXExflAjR2jjPZFHVLCpgvken6vxp4udXNbibLl/fKPrLSfphIo+FiGtuHTaAeee
x5ixv/yJ6tB2x5Xj3/oL7FnfUBsXoz1my1GsSni2Mcf/Ocdunzsei7QfYJ3fW5oaYZBRlSkldfqK
vF30c01pczm6M4CyGDFCr+OfIzRetC9BKOHjm4y8L4NBWg2cptX1JRGimpf+B6ana7wW7/RpCorg
LCF1x/PHy1BOa1oCyM3SgE0Bl/PeHHgSVPkyr+9dWSuMNQTNLRsYWKHceky5ofStCpbVfaGAsdg5
YXrb9GHALMMANdj8B/5SeuSIAQHtf1VngKBy0OxC7tmcmkDHLf21htFeFgliLl3eJHjPS5ZeMdsp
Y2q+i11YJmvj35uotbPhgVeSX/Ks2N4lKurAYebWZr81E4LLngozL1kqUwDoDnVjOUXnANNokK1p
p5Pl0mrop3LpdoDxzF9Uw8xXCqTOdUhRS6HzJgpjJuiDxbgtI0th3m55+BDEPctGhCbqVF1k6iqV
Gx8kFaAY5ZiZhNWZJuUH4F/DDn0BXCKzvmj4USlH89smB9sqW0MDzr9TRwhuL0AJNynwTsaYUz+M
ntBqr1kgoEMoCKiDWCv/avwkmo6KxCb9hg75t1BkpJGngV+IIGKApPpG01hO5cGcthkZM8Sg3nCY
WeZyewDK8MXEBRtEOhCG2OKcOpXcA7lTFcKgu8r6/YGnh6PJpd+j8kJEjW1Xm+0W7/r2XXSNGf/u
p0qSwClIgHC6Sn/5M0BCUsYtiI/X5otSCR3fumXes8n3GrKhGnhC9ayyc839KNVcHGsSW9dAGRoS
UDMV/SdTksmszAjSLiXK7j6RfEbnQEduXpJe3jPEpoaNg7Wk5m6yLeEYc7UBR6YTX5kTa+CZhEzE
ey7eUOPGhi2XWeJR1ohV4n21CCwRRYHiWwXsdUiAKK8m2JFOdTmwZ9dC3L7EygCLrlCefNrsIKpg
CB42M0874PxlYmvwvwLHWnXP3dt9yANQIQSl38Q52iLc64p0mkkkGyun/AoghqCzqL1I8PnnLaLI
v6xockBdA+oOafP/yBmBcyHveh2pJzew231DWZR6USOLUDGkFKojOrdHEx1k5VnKWl2aRTi9riBl
Kl6SFpdAigFY4ytRqp6BfsrfJp3RKfFJ0b+o/DmQo8rmFPmQauUhrW+FYTPERRfjtKxD1+6pUgKF
YXgZTIhyOtwecfL6GBWhsXCvlxvEyGo8UQvn3/n+Igz/8r0OPvbv9ad2xwH9YZdkYuRZFUj2p3RX
QRjzRtvyWmydVe/xAjqiZAmBITn19lmHfkJA+fUpETcGdVnviF+oOqdnQ5DEoVp0vkTcXnAwTE3q
xue5sVaX467OOhDSaQcMaIqSqoIjxKGRztt9fWj9Hse8ILQS7bfRIwqBQpJzEcJTeCtNdLGEeO8T
LGYrF+SPFYLiAaWstDVh+vhArV5FoDzj/dyjonI6sCRVL1sWnc8UvMHOZFdySsByA0B3aE/XTzqb
nGQy4KzzQG9K860I7sJxPcYtOu75QOuMUst4V6WnK8AuMtksw9a6jWx2BnljtH75042hyQ4Xl5Pp
AHRXxnJUzhwOArDZlX2n9uEajGMSiX+5GuDH3XnPG8jcvDM7NLQm3pa4MgcqQ9+wYS1c7awqki1D
C1vWBSq3m2v1E1bc1Q5Hw4YStBzcOcfKLdJ37//ZVWwNCy1/WXdERox6bYO/5+/9YdSsPfzV3dpR
gdQcrOKsBH/ngLOHVCXjIHSCvesW49lu6iPiOCPQowR3jjry10h4YlXPWiG1TKc0SU5TiihKuoKJ
Fbr1RGDin7VmQ5J0e9flWSzC9UN8HYbqzpKQi+cFnJJ27bTHno9cs+PRCPP7HXc9IfwNYigDIFU0
jlmYfjerSlbhoe8gYTXR9PL+s5s9lmxFSTJMDNmbgfd0oe1l8UCXrlF7Xyagwq9W7FRGL75t1BL3
3rJNSKN0zjeViKtuoMGQ0b+itb0SBEzhl1ck9eUcEDT5dQUDP5NCpHr9EK072eDYpt2k38rbeijc
TClN3AHfg1UVysGZMq77V9bJQ7IrBDkQUTqnn+29eM6g9CjlC0OT8BAZUCACLs3+RiOcTF7rboV2
BZ5zdDl2n3LWLDeWxyOXuHFTQH9Ysuko8lKc3xx6djcu1uJt5bYY5rPiRjlTe4iZ1kt53gag1vI2
Hw/I0h1bMIjNBJB8MHkNym4QVIhJb1OCoZuw1muWetLWsx1zP9hHCRFbq0Ku4TTfoyChok5Ja/Ox
2EtbHkzB35lWdWjwjuP2dRRaD23wAuUJyP5GvRfMjzP5MZHD7rHhr1G8XUSxV2amH+SrDsauxaRH
zJHXrKTGluSjBJd/dOu/vpsHksiVj553k2U11GrY/kqt+/oglvEsSlpZYYenrClMeL08zhGj4mgo
pHaXtb6YeEfk8p1rR3MFElZ7byHsydoi7RSfMzoLMGZMhtaWH8cUbM8eBXmHQjGPhvC9TO44zREo
gURauv0evjm38QBKdfVEN57khr489KUm8j90trZjo3u5VZOXERE1vD6D86NtDds9PPMqbjaPvccT
sMn/eERLEmWQ908QW/N7mq/zB9KTQbmjJaz/JBsur0LSA7Aw434JB04WFK/fZRy4S63d2xCsA0GM
1wGT+IxguaUeGkDp00rpmS9w7ZjLcmH0xpjHEyWG0J9/VrfdohC3GCEu7hj4WN0PX809a3E3Fq4s
ltF5QVodnaVr4vJAsjY5izdupYM3r77KAAq8BIOIPRxIq3yE0ZAwsYzRmy1sIhrV/YWPEGeAKUBa
K7RNh8ewB8ZV+KVJn51Dk9dOt0a9udaFDZ1xh4xX39XISb9xrE9UZvvkJ9JWNjEg1H/RH7S74kH5
mw9nx/MFk+xBZf92uS7YnvrhlxwU34q8oqQJPiTNrFTUhVCRmz6mxq46Klb/79q0dlhDGsHuMXB3
KfMbb/y4M0FuUicJ1jZRsrKetMHZ5f4BeqR+OZ0s+euK65czbe1KUkE02Oipmvg905fZg0mozWmq
PaTN0rEnjlkBdOH4qMAXatHvZs1c4+T+Py+K40GQrpxuOKLZvUQNODPCsB7DW8Qf9Y+EQTyZ2xPy
MEd9eTDzDGqhZCCZaECbgvDegC1FT7g/+CpgEpldspXU2fZeS6Rc6KjJArXrnCBcv/Emxx1qUeEP
MSBqLqgvlqeZEttFknwHqr+ejvkW7yiB6qQdyjb2bcf4PHpA+85lm3TDonWAef8fzoU7bX7gN5H3
AOs1eQQ8HNOphdzYsJhXHVZTPxHo3UVqVPG38J+gRi/sPX2Tzhit7R5Nr29F94Vho55RlnkzjVt7
DzD5fbAD8GIuYTaTmQgxf/Xhay4R/YKsnJKo+NmdO4NfF/hYoiLhYJ0s7SYr64/Wt3qAN9ChPY6F
d0VBLQy+svJnar4wVvZWAE2IE9Do03qtJC+lucPxDJtnTcwGYXI+vkn1vbpvHWAUShwocP+3tSpH
+E0HtggbPlscTLsdvyhJEwUeVT77SbNgzFyicSkhOHPU63UA5rsw/bcWJpqiofeY6BdDjVpA6yZ0
39DbRLp1TIXTOx2j3eADLgPHrTrp3HnaYNBnPNDcIJcMfPoZXAsfVLJgOzulE26OHcY7tkHzN+OM
p3pReUAs9ODuXeuR/c+GcThEEKWDMZlIit7JuKFYieXvVDUdHJR7Gh25KGCGkcA5U4Vy77QR2PF+
0Mv03X7yncrWbX7sEr1RMbn9RwX7orbMV4CM74gfIa5vMufdPPaQ0vM4qw/TpFdTwKj7IUIMUiCA
l4mehsnFAK5gc31wSEZy/lcFz6GLu3wtJvzvETQStn8mhnbt3DPm3K5VpKAbD4pGwVJB2578yn8c
zQs8g2oYjRHX4vs/rQfkg5hNeYz+5kbau5zzvd99
`protect end_protected
