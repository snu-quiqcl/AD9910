`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BQ+trpakb2k+k7/18znq0wwe1zgXP+hUt/IqwfZTp/lGOe3COOcIN1ANJOre3KaalIg7J4T53q2y
iIg1ahfqqg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xXnnDpO4eL72ohheMotYmgsm7YwJKQT37JTIATPPekNvaNa/110YalIhG6eb52hBvSDLJzwtAtzV
E3dwpFIBZJIYMAHzJTvbhkfqLD7/4pPAPBHhZQNyQqL+YbC9o5ydTFiRkWfXAlvJymAmKAoiIlTX
WDYEEFqnJwGh54z6e78=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FkcfD6AdnMzzDK+dPfRQM6XxgT5RLRDECxjrRbJh9BV9xIFXPLkNYL5NnhW3ojyIRqKnhBtFTlaI
qtaBnJ7VN81BRTCLLBxB2Nzm/sdqBG71nWZlRVcpRbHn12SLWbkKCTcXw8jDE+JF0ILLr6Jp6leL
LR1TgAMRa7y+SFvmEPPnztSPSJEitTaOiLvMO8HfPzEA/IKZ/Q/1moLX99mxOVpGVLokhxH6V4WD
y5h4tHArLy5NSISeqWJQqhQXIddKGLiYd5jvh1AAN6jGlXcWCCxXLHljbzmcjGTpKHUVnGJ+iiTP
VFkevOen8Ryvn8YIbzdG2+ExvKFJf3cSeMTChQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UIjONl4yYzxEsi6/0iyZbn//KWstHMZLnCjGBfews6oK5XBfORO9WiMfxyVzxg1wS4ER2RMkio41
Wc6hAcdkZK+M0+gCWJmeqQj4Ml1mGOFENJKyEveG3J2h4LoAhs4kD7+s7kPZOZsIcFgZIjnoGTlj
8Dgg0mSWd9Bp2rBJ3T9vg9QJVs0dbXzP7qS3n/aX5+Oo0I5GDYl8R+jE3OCCgSBcUrH0fhyKS53k
P8CRNgtNSBqoWoewlyStUjundqvchV/ZbYqvjGSqsRX3yoalOyuFqmHTrNnZy7npNFdZcqqdWshh
3sODyPjkhAmBHjNEx3IkVMW8DEenrILStXERzQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e0Wl6FUWxyprVs/DoAfSfBLzxfeowNuF8hUuqlr2IZa5Cz2OzwxmYBxLaFQg6ptgByBJZDRzup1X
U60jAN/Ug5G8BFT/jL1Mz//awFyj3EYnQ2fTt/fojCxJbaOYDz/jj4KM9dCPRMYpg+MHHhtzcjbs
VYtryZzg/zyDTyFcDGUp4riElLwxZgA5eziwR6UfbrVyvUcuN8xcfxrvjRr3M8wzypvPhrA2I5TF
Nt9KgaAVzSo/YWWxoRRLOVEPlzXyIzpxGMNMoURZTuKy1lFxMsyZmO2O63lEuYEicNVL7NBt1/qI
LiFgMgmhI0Gh9B8QbBtEZS4bgCNS9D1lifvSaA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G6WPln3uw8TMTjM4Kfa8nWUixjX/jcnGVJqIBJkwcRc3HLOduaxsWjrgipgjB7/3xQCY/zpIPWlU
yx81N1Eqane7gIO4xHGGUYJ4TnTZxVXkeM1ET1i8VOvFCVwC8n5F+n1kLIl0gU66YgrUU+LtXHHc
uOvP7viCAi9udgthQ4k=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LJ8bKEvLt2ZZ8DOv2510y5MZx8di3DP2iit2iYL+j3SmVFb4qDP3oLwF2iXpxssRtY/FH+a8vEXa
qHq3HCl8F0MUjvG6XGlYbeAaKEUiLKqlzoedeN9MjGcR3kT3unliIk3qxmAjmcDBeErfly3WSUmJ
N0xd1OhDl6j5F8sBseE41abu0LaJQtcCvUOO6wQ+yvyWmqHXOWDHjvL7/lLaloeCYWDrNyZDRjux
ZDjCzEvudUUS//TFihJjAVcuHw8W1oejT+HAsJzI7rugztkdNYonVZid/ThjaBMqTP0p/3naEoAt
uIFv/JuUKQGcPzWgnI1aEuc2VpsGMWQD6EGlLA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121856)
`protect data_block
i0CDZkMNv5O7kMpivWDEnbMWZuvmx3B06haCcdcWUe7LVWiKgYliPUc+YkCAocKsqcW05vCkeU2R
MH7nQG8Ye6pkjIlnvlu6BQNHUpfTi4nahxyQaQJhvHj98vgB7skWz2wjNyhoaGR/1BDWABwNu5j4
y684CUQyQuCPhdHOxksch+HEkr2HTbLEpZStb54cwp0R8w0EfCkjPL36x/nz1VOyser61rR/R/wq
wncAL8NYKuxL0NUIcQCz2m99+MFaw5q1cl4TNKR90UP+bvgteVxrgyINXdctWylWP7HwHHf229MK
GzLknnEa70VjQoonlI/quT4lcr3+dba0gOWI68Jx1m/8Xl2T7of2C0X3txgLmpBYah2/WWerKnrc
TK54e3a1i9v93P0KvkJgOy9ojKy28Nc8NrzIGpvUoHozLUS3steac/pwdmXCvtD1OXfsfCCySQfU
9IfEntkB34RAy0qbtRoGFZybvrHVGSu4AZ17raOiWQStmExxL9CqnHdmxBQXYfGqe09xstCLSm2W
CJsk/ijPbzMAPh3Vi1n/3D/bSEL6kSh1i6lpzBruwZs5fCooeesUgfAmhma0DNw8Y7INzDm8lseu
/Bc1h2B6VcuEuZp5NBK4238OkJdEfrpS9rznvE8DCOrrJdglbBcGzIc5O/RJTADQ0loVGhcyKALe
WRp0Ha0S7NINyc8/au3LWEHv40a5bHPvDu3l9tRAyXUqMeUmjqDcI1ybWfWKJBLVx9hrQbBNM0l0
E881VnETCIO5lxo15A03SPC03lJHe9TPLWJJNZS4WCaYz9istadabs35DYZVvNLblc9I8eUA3lhz
jRVEH272Zrx6uVM63DnTiCJ/WUsGCBIRfDqhngJ36JHmL7sfT4TLTa9yA3ruX9ZyKCV7n4uwZ6Ph
/rcpUv7SM4VIte+/xcvsYr5VAFShwrZ6YfLLN+N23Is7a9YAzdRDLJBHsPMM9r9Z55i6IC23WY/Q
J6MO0mKBI9uHy/wgyCPcabTWKYse5WwRmnVojNgRCuRkrKIvaw1Hn9IGjEdxitHaTUIcyXMACLrB
jCmRRscEgx/RZrx34dh3li7+CH+N09UYuMS8pXkKLx4DTerAPJmXymg6tzkgyR23jMcPLLTsX+FC
ilhNdx5Jm25QEt3+/alu2l7NLIUz7xXfk9PbwM5v4PFyRLCASCvtiE0dM+nV1qAWIwNglMmOAKI3
v/u4b/FuPiR4auPYEm5EsE14ZcUgnD6mwDwGQSXj61ttuzbspqG9vv5UItjffxipVyZpNqO03msA
tXgySOkTrc784fNpBvtQbQqwXIR0oLtSXwWxjVz4QzJJeYc5EO6d+Czf2VB221dDFb1+ZQjVdXCk
BPokUiWX8w0RCjYGV6LjHCeCmovDYTXOYRx2ke/fAbGFZAPMyYFzj1Uuuj99U1tk+Vk/w5EBVG/4
hmQ5OtLWPk5MWz7Kko+JLoiEEwp9g+jJEFqHGzLdqshYJaoDkcBxtG8wHGE6aLeRDxTz1Ewmg3dr
b9Xmu7KZohdm5h6a/dMbWm1Q5/DJBxQUHg0WOF3inHxfjTdger7PceV7oV0RtypT+AHFx68ou16B
M8tuHYjMGOw7htE96jt77JdrOXV86Z+ZyLUbRJdXv3mA0cRKuCX1rzjuOv5qdxR7XzCcYRjekL0o
TFL/JPIGpJed2kBS7iCqCG8Iw6xbAZpUJ2Q3nH+71STdwvmVVTJ6nJP0jzxxQsZh1xZoY6M4KM76
qlS2H14YCbu7TMT7Evipe+9VdNqVc/LwRcxev/Z54l2aiVnjE0FKAZ4zJL17dNYBWKkYGln3P8yb
EL8Guf28/4fiUM8TBWQ1zP+LhWRH61JxeuTU4OlUrSV25HOdwg4/ln1wl4mQ5WThU8cbxxvqQcUX
2/dmIBjum+sWMwdox2hxo4u6BHyjihLD2JVPdP1OUW3dbFf9CVOoS8quuFR7KDEUt2xOW0388//g
6VX40M4o5LwSRwPY6VyNVthZhTJ2QprQlxf6LLo5poejnwWTAa948xE1DDfwtHB7Rk8E0drO52oN
8ffpVETiOuTUdACuhKlFXWQ7XG77hUVjxNCr7M5N8HabWL+3EdBvAEXI+btzDbv7vNauLRmWGq8w
rlyhdYGZZqcQHWl8H4ykUwE+xMevA9lyMS6sD9/bOtUNsI8N4oxEb1BY12kd4NDHTqhT4FYekGZ6
8Wv/ds0BNOPK1dURThUsUxJOst+X4chDsMVi58gEy3Et3CrxNxmyZYV1RgL/mRe2NxO8q9qYxKvS
WFnMPeOCMa3nntXo0s8ZH/Y0Zla5+bdymc4IxRYDCYQM8MBnWg9KV09QtXWYIdDV7uxACktarKIR
WF07wtx3PEmSVb9O+8AlKxCmnr0onWZ1isF4/xagD2Pf3n4ZFlX7ORhA8kuWheD+IY0ZLkrxf+eL
c0XuyjMxhuQuQ5cTgZgh2SKBEWaTixKZCIqZ0HQqUx/JplbBHZEUt2uUWbXkrUJiTwjdqd6E461G
EnSHzIl8l14yp03xe46md8+pkKaFV6D/e9XgTShUqvVdq4WTvgyLnmsU/et8GYmcIePK3WDdDESk
pQz8d5EvgswRy7n1meTi9xueB0nTFzlsed2cWNzjVzYPNFqgrclelgpUL3kti2LsnhQH4yq5w23n
k5+zHhTKwcYazTxIby4vCz/jPTyPDRsgfc+7EXiLD11wISW4Oqzmhz8VQToZGTCRChJRpqWnCcji
0ONl7oQvhC3dJZ8yUDn2JlOM3BzmdDwW6pkJ0z2N5dD6ypcrHSN4DyyMjnuND9zN7COpmL8HS2Qt
Tz5kx3OdDPYn0NCSH00KUswODU6lS5imdaZUT6xekdyDPm/d6dccHnJcoRLBDuIrEis/CjgaJRBD
Il/mWnazONhxejuhcjtThlvDbMY0l1ZH8k64cxm+DwcIBLvLLCY21emKPy8U53CCLWEaQDLFOcSM
hehsqQDcdbQ98P9CZ44NvOOcmqqTWoBUtgQf1sHta2+8RMWH4QCKS5OBpivsEno9knkqt3Tygkia
U3Efbco1ZeaoauUkWLF8k8MMkkUrHZsdt+JsAULhR3X9Oehn+N7IoLQ1DN0RVEY3wNU6hQBeQSXR
8WmznsYWVFmgkUEiDDRdzVVxIFGHj+gXzZZse3ZGpGQV7Sw/HacKK5jMfaW9E2Uqpyl8acxBy/pZ
c/LuK6iUrFoqZVVN7rmd+IWvexe/n76fmDZYkh546JbtXmEk+ehyZSm4DV0jZkIe64GDxBe8qEjd
EDKmEbOMcEZAug3PTF55VG5hHofe6h5+NMnPtKw42+LfpS/s69AA2lZ6glbsxdLZ0BnE01HDXLt/
2CiqFYQd6boCYDc/3AlA90u88Nhtmz6H9VhNPZiPZEnQjpqwBHZ7h5HYz4co77i9YCcdpZiMiaYC
/8P0KBgGCCRw24wFBuGDopIIrOCV+BSe1jSbclLdt4uNMkLA3+90HI9PhTk9MlAlFku08i28PtLR
cGnt0a7PZY5SPA2vrwtAUjvtjqcnsmw+5j4neZZVJBxaCOjSJuqbao4MJ4c9k8nfPYyANpS8zh5A
i3qaNhQpKuPhs4elktk4hVwK7MMUYwAIahLn+9FzxgTRXzkYCiDgeX57Th5I25vt1qq7GWtOzN99
147vBcgDFfFg0K1H/rufQt/VE0TGfJD+3e1o3NPM1DPPDS1nsone8JaG2o165cgIYaDxN0GAiKzH
oGPCuKhDGxr53rZvK0PPcvfW4OyVPF2H+ajxWNAveSNvl8tgLGAb10gu4bvGUh8dL/YLxwyh49Nh
iTRm+M0GjFWk65o+3PCzmhpKIpv07/JH1PHtfFlvxD44TS6pNsJCYhQsOCyZP2pkaSrYicHngDQH
C8tuafg422hGmwhc6/Nxgbyjysb7Z2tMOVhSLtOrSZY+PKBToYDZHWhcVnR27oBHdjyXqQGPYs5F
PPS/WlaxkHQeQWhj4XxSsLju9imfkqqY8NSHms1mBBEH15OGv8QQoRxT5O3dPNxEXsRGm3PBbFj4
KGykJlAt5nNtxbk7hgqIiIFw79q7DKwqX1luVpwZRsj8oaoQW8KZxNJw60UMBoEDLrtrQ4Gqc5s7
YoJFOBwIJvA++AFoDuJoVlEKJsT7glsKZ0sSduFXBOkHO3LZsE+pd2O0q3t+BwlO0jNnUthB93e5
QIfz6xXjkm/ZQvs5PNyzQos7gSG+ZDCwoLghm/ez/k+/yMuLGo+P//B3PUjmkzzHhs4RlAbCigDK
MIhc3aO0qx7hS2mSG8rBHJwjBMvuPG0T9Drm/UZWV0VAVpE8ex3jQ9xq4i3fotbrW7tR1EAp7RjI
c6IHEQmLsw9+S0J9iD3AatooroI2jgyK5vJIYAkAxvx9zxFNVvIoC/1JO83nSZQ2taWZM4EpjI4Y
evgBCozV7TNrjPLvM+PvwmsAZpuvDoVNLBEfxMz6L7Nr30hferVmGOLeTdSLW7iVKmTIn4cEH4uY
j7OOq5dtzK1OMmDk7yXx0yb7ZWWLDhzgh0YWRI/1pQQn+c6UtlyMBbxKSM9ElM28//9rEGnTyaVX
XuBFkzd4isjDeKwgBeKKW4YoSRN15T//AokNLF0VPxm3u4fluOhDfdUKVwkiLPwPtX1iSh1a/cM/
D4LoizAQ5BdrWGDKmDQuxSdqBgbI665dDlkqlw9WyJ4WnBKN/l1Qg/HM5/olYI6/ciU2DbXnWkAp
0PxcbtvtTqnndX7G1RAd+Awpq5k8xlKVsEpZjwFoC+gEO3NbwAUP4APC365DzHxSJ38HZ63TT3TL
Y7/N/cRrF9Oh94HcBOlcVTpLzO5Na1uVNINbvw3p9wwiJ1QCOwEieA/W9L584EcsVY13FHUQrX5C
Ins6bn4akCFQlYWYOjei7ud8aNd9lj2sUuclUTiH1Jb04USm3MyJgsxyv/HGAmmnr2/JfRzjp9Zn
KZW9qNDW0wY3nFzkVQG/T7+dHVvVkYb93YE16XzeMPuRR+h2gb4ms9xWwxCldgHtXWigvQFYHTqX
esubHoq/vbF0zK9kSz0Ph9cib4fummnnFAEpydInS52anUYNMMnIv+QP2gBEpSj9T3lGXbWik9tV
3yperKkjUW66JiqZmPNyBRlewo+m5tFDNjwqB9Ut4PV/48fR0apIYSR3EOKfo3CzmQtu0CEOVkCj
cHdz49gCvbBu2EjoNliIZcLXfRfElbhKpkHW/8T4GwWUzgIAO/emtil3hEqWues5gbgphAmsoo4i
uL77Pp575QToPp3cF/soD4bh2pZsKgFnj2CgrhcTp2arJrragMR7FSlfm76i7gfUA1pVCSOGsBj5
nidKaXd8XcHzHo4h9UfO5qnu3KbKFa0h77D7CPahYE3UlfnoVpzsjo9KcGsnMoezNP3brJjn5jRj
XEKyZNeHB2lHynvg07AhByn77KUMLhiIBS8lwFQNaurfURgxOka/g7mj1Jaqz9GqQVzb2Ic2Vs8e
s7uQWZwnQ9QC+82Yw7UngJTtDpTO8N26GGmvOHZ5doskKsFSr1bsNBuj0MjkPutHLbpyJjJKoydh
RUTp2FDLaenm5mW/CaISE3Eiucxo/BA2jjCQTzVOcTFsMA1gMRaZj3Fpa8WESuBjW7fm8fpkFyZ0
VxZlGcrZZp97VJo2UvIN3kpCOn6LpYsxYUQzw8fspgc59l1RAFlOv+yBIBcbCQzBQLsNByTlwUab
t7OgFw1nY/o2LJBP24eGzxgfmUnY25nnAgQPXNFKnIXBUarJXqxHFDExBk4dvOAvVslEnAYaP/Z9
k+V9cVu4VwoMg6VAvy9HgKeOjc1uIu8IZUyQeX/3nqDlgClzX/DsVRmTrmnf/6TR34UU04HPsJiF
AyGND0xELZlbHzw6yNzazqDUM23PxcAGrlzWwVT4AdJhlcN3m6lhLMsnm4z8K9Oex0D67CYXWG5c
lPmDDdOUFko0oXe17nEQebQ/sRVvuyJEi2JUFL+oyIHokNr+r5bMq454hf0OrdY/RVtRxTp7uPNO
DGFsLI70iYJMRdYNJMyODj3qB7khp/9FSG/Aqwhzn3TC17X8O+Q9g0TLV5ltyxsg/9oaye2LGPHS
LjIU8p9NyevPk/0SQq7q4/eGgcYG6CDPOnvBF8fZgYlSxecmBlG8f4Ih+eJuas9xlW2LoF4kT+lX
LDc0oGfn/DntcASXMPtGcMoWE2UJ5T9G2WtR5qBob3nuijR8bt+r78Sr2t3N8tLdB7LSSfCn45OX
0DsZXCQ92dKXXoyKUgG3OnpAKLyzDAGXCp/JSl+PIGWcfbqkyhtfARXd19XX9kAtjMFespF64nvL
rZs76B+I2QWp88LVnY08VkoPrkVoaXmmhRquGHnjsfxximrczkuMdNJgYj1uk9u5qIj5qRJOR5eY
JlC6SAE3LRT9TtJKQTv4R45qnuiAkZOOUWuHbw5gcTFEHjWz6zqxicPsy/9Q1D7r0xqu1q9zlrAO
Ze948kJqRjr0z/O893ix2x7PuRMQMpl8UNbbD5XDJGmbC8v+c2JTAk//9EfaYJ141Pa+7W3O3YnW
j45aOH0yCz4svH/R6E5ORrQosMPD0Lz4K9EKhRKyBPggqkkNom5xiLxEM2V7XIaS5Cw1hXVUkcmD
OSlzTHlnVXjOLSWU3NN1GmSkH3etHRq9gTlRwmjKu0af2IxkU41x+aamtM0h/uWq6ClGS4jqPNog
P7re5answVqa40kaHN99ToobB1lMffNR/gvvoL9E2EBIzXEmcfmmxY2wMzwqwsKIh4+QdoyEvtVT
aFN75PHPGUu3jrpMjTJQ3LvLKA3jxQ2ZzQPudVJDVTs4RhYIb2ffsLpNm+XFOerMlOSA7oOzcOMM
YLLBK0+dEYQvyCBzrFsb6QcOHQXk1QIV0UrCIayHeVHROD+O9XgLOsy4HL08aFuNaA9xqbYKtZX+
2Rw0kZg7i3ZUz2ZCKsIim3WNAEdytq6v4STeubO46Jpg5rWBKLvLURdjQcyeCQ9Uh3BPSaJAc8Fk
t1R6zuNd9UY6/VRG4ZhBoKfKEN+WlxS5CYiUcix9Wwn0I0+MLCQAaKOGjplYvQteZBsY7H0D+5Mx
SPI4sxPs/HCH1QyFEP5TNZ8Mp1RlczLTBPY/0vNUknV0fsAm7uSGz9yGP6oR0iP6herfS6qQF7Rf
zFkPbV+9Igy1wZMlbjA/RBLJoP/sxZ7fZHaRY4cMIsWH0gTradPf77BsSlTSTMyd8gRQqJzEyV9A
zblIyrFILtaAHPVSjhQSOwOAciqm8H6tMzBnprFwP68xJpckw6wkk4fR0I4PJ2EweDaJ/UUFTTpz
URwCCp0vpVZ45G7yGS+iK3hDv40z5y9QHjXY7VNZTCBTxAN+mkGBgPny7JVMbYbN7Ez+hgamVK4y
h/Hqk9cGiD8azhEPfoyALvKMk127rWx7OxnXQKNeg/5KvIIfdxchXP39EvlnRH17i9q9O6vldSg/
ZNo53orkrOCRpJhZ0adcC2MW2wz0WQ0jl3aBb9s1+IOj1tOMPD93jn5ffUaZxRlfljTUYyes828S
8tRNex9Cq+CCveErw1z8inpm+sypKsrzclHa3n88Ww38V4i17dS5D5IIKdbKfrcLbAwSzh5VH7Fr
UvK6L6wzBASE1ylJ6DtEiz8l9MXgMAOmoX9y5r329GEh/nmrBGTVN/ZjuWiRYvPJ80mPYv4tTtHM
fKb31hmE8G13Mi7iXNpoGt8Ve67p9BNQ/p5Y0cJ3RdZ3jpZJiVdyr0hnNknUwbV71rvcV7sdQuPR
lSOh6E7I7i7bBC4oCXrDgyBI1rlKJRvc9ymeacU568o/4U1jXLqO5wLxZ7ufmCj7KHPURaqH9qUi
8lC17WikEaoq6Dcsv5D5rvtoh2qNw8OrKhs/CfmSYxCjHqDK1CY+ctRpgUAYHj5elvxvCiIuU4j7
zzeFH5o+50/1tPMoKgWfLdr1yVTo8ziOblNC1hefB+xovRH6BBh6fjH+oEVfEAYtfYVZFs9LOOcv
dOSYaAXSHwyrrZtsfdCdHF7dzGD3PazJgh1NiVHQFcDDW8LbkoZQPcd8Ee4AgPMVEpdaFAkD2JiQ
o8d1DP6Tqg+v9tiHTMk3Ll7hIUogmLJyfVrSnEYslKMpvZONYv9LUs9+FzVV6myGv+3oPAvMzexH
85yzObyTH0CQVyh5JX3xzyTwRTE9rn+WScDqarK0+h+9At9RMXYxEBLJyHJWmd4zuDIK9qSMsumI
u//6uY5czTdbEUgI0HHA0wfU1tLwbQmApA0H67MbKoQRrJgkZ87Ks/c48+7llfTA92kwxi707lAG
KzvmJovcbuKf73YQaPuWgLB1TtdRXDz1HeE+szgqA3Y5ko0oln7zlleak9s3rqKOpVZwNQk1Ho6A
zb4od65Rv4NrYhF/99yv/sFb3zFOL4+VhdjxVuhwMkfHh4on56NPDkKqV+rt7oL2hXl4zPz10wrQ
DJiQOev9kFw/n4tM7j6OhyBxZEI9fpg+4kaaJquii6gcLvwAhjcK469pvduoTeenrTkXGrvsM/MD
bOyhYazk1NYUOwMCBBRlDFIBao5EI5y47/KsOHAx0RwiGFMCmRECbidTpo6heenH/j2p1/driIV7
9t1e0uJlV6c6QXVfAoS0/WuF3LpgDgQTZExEOiGTNB7/CSZz8toUqF7RR0MsDMXgDq9NgqA6kpWN
ha+yMqCGaFboZCEhMrv8A7LOSZHWsg2CiGnU5BdbWXvuq6PKK7xnJ5AR9EkuQif7TqQzJhiRQeHk
xyGHTbBSrw8sWIz5owyHE+2pa2DEsQYsXdNGy3uc8Hax1/j0hSX5hIy34g3OpWG1755lr8O7hfQj
6uh9zkO2lqkz5SZL9472hhPTd/uJomFG9OBgGTNPmjcAnlWkjVksG3G3C8oaqImr12Agxp5n0UB3
hZhgD6yla2Fjp3zmcMEmy0/pRBMo/KJXenS/huhxTmWqrC879fAoJ85LvfZYqoEJoaMWzH30U32D
ZaMe3wATOAu9JsrUmYbKrSNKTZtiyMqghf4t0Gpeg0Yi2mPyyGPOwHCghLHH9YvSDwsE+6UbZ8YV
xT/LlZg8go3lYgKpHfJEzwG6d/NkVUqI9Li5Smj6lsNghuzZFc/sAp4HyWWO8cCEGwOkKn7K6hIi
0K846LahHPZkQpaF/iB4ajWb6+KNQSyDEi8BRTgmMpY9rV5o0Pzz+uNgnGdOtyACbWe0qGVMdj46
sY/+MFbiw2rualefkL10NgLCmquzO3Sgy0fuwcWWwmUkpp3DIBNLY28+J/nsAIDiXWAD7s1haQSH
ZQiz4sIJO/MCzPpqa0eShpti1ZG+6RdHcVTVYxSq4cw48Zv7ZfcKQX129HArpKRjclm9sBx0GmLk
Ji6m1DhLIiRh0BSxRoJ+sJHmZESZfR0G+ugi0LGnVKik1lLk/DcrenJIl07ffY/5EOUwdEb6Osgl
iqWXhJMxr/sWL5/oB734W26apITIsgIdUHJWAgSSNWlUQjBbbgxeuItRm8M9ZrzjxGTetZ61rAA8
oxYkXHo2haElqHzhGGtqD0xNXEMrlABuZFSJ+o7wlx7FHVcN1LoZ7E+pZydRxMT+uG5sgMxPU9s8
JdV20zmGJRT+1BNqA+hMOntw5m7PuCdPF7hmIXfHKuuBk4vlXQjTIA0/O2xHcMN09NT2xpLjsnM5
2MuR06q9y9rYfoMMU9H0jwCuaxB+YzuDdVKmwTJWfeQBblp9DwKlM4jH9Asb/je7u2yetleVLlIz
tb1Jdw73tF58SNt8FuJPPOV+btA1allC9iMDazF/VzY3t4BTgzy+vh2QCV4TivLcVEumREdfMsPR
DS6oRjksoEW6zpGhf5crCnLq/+bvtI/v9t6PwstIxRqkGLLpJCpexxmKusYGIBGJjKfBWB3SANBP
Nz0m+JjRYtiDf7pAMTVFILpB9U9KJ4PAvvQJ8IMxAjdtvSrxA6gLKO4uvdl+fjjDvm5fVcqiV3OE
F/qV8BgcyVLf2MU1nfDaHD70fPH3wcChfN/bnkEYf/6oUxpakYLuOk5j+8yBDW3mwFwBtlDgsZ9C
B2Ixc6L/JHS09nPGkRCssi7qDe14C7xhO1rC5bhnWe5p/kA4ZhrXgtYzONiO7yLv4Z7+++AmWU47
luy+xM8hgD66Zw0xCoCT/2ExnrHC1WsArpEiaFix/RbRtMMjrqeLyadMuSDrdL5/3C0Q2PiJhv1I
Jz7WckvSdzmwhI6d7e94URBtRFubG0sUxqN0Uh8LPWKfsAJ2t5JJgTJY3rZ/MIFr6IFJSFJT18r+
0p1CjJtNaTncbgE3Qliggog5feSWTnbicX71zcCYKVTNnEMxYmeNCVcFN/ZkyeugGFI7hY5GwfRy
QTU6yf2cJyMCBHXxNi7uc7XdaQQLLypt0WvXSpIBDVV+NuJFQXGUewLhEYDtcROx0rFr4Evu4+fB
j1tb79s4bF7mUdShcIRpstJG4JLMnCVrK2XGBnytJ4f8TE5S1xVRf/dlbdKV1aj8iApGlty7oLPW
zrEwq3rn9AiAwJcHxQNiBfvsrq3zpr+UUCCV5KYLBGta+dBQeGnWvE3I9JmlPWC88H/FBeOXTa7R
o6vBEhfFPKUiYUR2fl1UDano9l42+DWd3usgc5dSRzo3h3P54Dpbl9dB83BSgbVYFLhjA30UV+O5
JhhQOjE2I6jRnCTFKzpQ2yn4ic6IQeDWaPLNldWi8S6fT4RDIESdfL8/5lVXzbmjAx4LlWGMblFt
fydgesPJ94TGAQEGprZe9dYwU6qKtruislnIvpHl6A60vVFCf96mM845DSOow5j2yU1Xy5M13Gdy
yW0zLHjo9WAQHforF/ToCRU3xrErgIpaxzcdwyUep2pztvqe5M5xGvmk3eT/oKh1a065dMFjVLkk
ZBTco0OtdR079TQ/lX2qKSDuiXDp3ESMHxaPbAtjGYNo4GAyzIGXSMivVuO+Iu1+xUstL3GATI2z
xGbzT8iykYXnZUanVDQfHvfbHEFJ1pLvT/LIGMU7gH9CRz49srLMP8OwE9W+Wu3F2y4JIDzUv1IY
lr+NgSB3PeyYyh94r4JE2uX1ru3Aw3BOJPKe+PwzcP92SxXwAbRdHvEREDdIQHSV9QaKagXTwjxe
oYaWI9JZk4zip56xJXvxoTilvLo2nzWcO8VvhRQ47jfPNTKcZ1KCFGgw49qEvm6zwRPqqVMuFBXo
wyegerWvBZ765l0q5O/WIUXQ0PLkPgrwH1JENKfcQFLJ/i/4QB4OI7oFrZgDSJCYEr9dJ4HoVJJV
RWfmLbY5sOsRtyFvFxLcEcHe7JJFAnCela3ROrUmvWQpJscX9uXbisSCE0IVOgJwTws+SRbszczr
QMzjdW9Pc8Pe2s2SV/+LhxFdEd++k0C1LIHQqVPAuEtWRcTsVBOmV4MWtvKvnjxXQyiWJ5Yf5Uws
lpSuHcdreqtb6RK1dCG3R7zJzrCtjpSlFn0NslaN6yOeHKAD26IKumQHN1qrhwdzOn7ikAjOackW
cgYptcwyaJbtGfzvNhu5yN2glhg3Ks+4Ym3MkZ2eFt6koV5EE15ohOPF4wHt8pZkEbkL2mDwBXq+
qGKDW4OCQU4ISAXnHYb6eV0GcuE5L3wK1z5+38/xaXJbYgmlCZzC0mxemvoA1AWebrOP/LXKBbxh
yHskyr+gQSdINpCqjwz/AKkSvmqNt9gX5+q9EQUkPFraRdTUPgy9tX2+3WEfM8NuZgroJKUoWN4V
aBgCViR9mpKOVLroI8WRingBMNOo1ojTUyjub+gqJ8UisyZEgoKsheeylwhWKSTPmrzWdXD9KR2N
vlKW2FsILIxhfHv9nzefXxTOGZvj6f/vLeWvo0eXezMrEAve3EoGVNFMo9FDHEO0042DPw3R8ea+
3R68ouJeNhSfBISME6xo6bcQcek19AX0wwCOT3Ye6b7qehDCwSfcmLTDnah9xb0yBcsOcggtBKxF
4Yb5a5gkzvBICkujqKir6w2W6JUQar76QF3fJZ/b5Gtpa3b7gnIgJpz+GuCD8j+XKiXBwI6apxAZ
uKec+L8Fsr13Tiy6QNLYhQ8ZkRThTz+Uw78pNNbMZlMUuoemKimRmOhSc8hirdQMg0HY4lNCcurQ
BcgW+Cnn0pjHU5nsWYldFhG1gXOtqriPE/bbbpiSSpuU13uWaA905RBToqbsOKRJh6m9BCdLCEd9
tkCgLoAhq3Dq8A6Bd8bB4OYPsFR6LY+cCw+pftXCFuw30OKpkBGJcU1tnmTAKCsfJLkwx0V1O9NI
Szr5G1G9lE8GXJYcilfDaZ2ytR2rffNQEJBP48qxdC5K9WEAqlWG/gs+G8zHIEymaN4grUg2sXpK
norhhh9mhMYVFKkKg01EhA36+cjUKihIo0++ufX3GSHdmF4hnKXFDDfoMi5CcKr7wsLgY7pfFbm8
cLtBlCuWnxWR9L9r3A1JffFjIMKMicTXf+ZZNWTftF4l4EqSopSRRduC+QzuOgMhbbGS4UBQd92P
HCvDa2CyZ3fpDMxiYPmsvK2pAL19rSBFX64hT+oT8pRAes8PlTGP9j3GUhiTvwXx+j4Q2LOc6+Bx
tlqh7M/1/ZPxPIUv83qLPaExj022dGfybgMZ/8TSX2xg8Lk1HLNZ3Xn3UnVjgRCOUlDKjarVINxZ
QoEZgBAzMec9S7ddYL6D212XE/R2hV18MdLAp9ZxGOQr5lUiOKd+QrE2ddc+wHbg09skCTBHaYsx
uESet9yBBa5tt+FxrL3FS/e+2FhHjebyVbFw8cKzvWgBmZnmlruNU91Xvr2htqCJWr1Z0C4/Eu7b
adwmotDAkdUA0t52cC8cgTXd2Mz8xSG7LtGz51oRmbVT2naesAPf1LTmnnIdeEvdC1/Yy/fUurIK
qzagNNqyCfmljp7pYjycFW5i9OquwyX22lobbXixlKKofTjUnMQkYZUFCblyTKBFOTtv0JgGTX8P
GOQo2y8CpeOK71p5Z7c4t/Vxozw2netuacQYy1pwT9EJr/LhZ9DqFcUWs3E1SDab3IQ6126UbVVc
3O3ua5OPsip6E1NVutUhKBovKSM7z4B/DD6A0kzyuHjuR/QIX4MycT5ycUnS1uemt4Uj73402ZlC
sl1bc5s/9kp9/awv42wGxwr3s8Y6r0Z/4r2VQBR4k6z/o9nrkAT8JRDQJvY4ubXDxhpHxtFbqGkX
/myZYfuNqQoJFx95B4h39xS4c5ADoQBbf4+l1Eoj3UhSxtGBKF1rKhM8S0hDKIRjM6xN75NJ+p9m
rXD6NbAE0dGmLDrtUcI2jZhVLWOWY1V+09emsRzXa6LmUWaeHTcqF9IAkMD7Wayg0A219SwkGto/
cql/npbtocPq5HbY012NdKDzDz1PVuxEtNONw21GLXUuZcoV2A5osDP8YfC+k9exXzjOdJwy/noc
ZSWMa5IiRMLB/s+OoCRaryKA2Ux3+Ic7be1Lb2swZWBBGiqvBz/KJXkfRxbNJSqyBoliaO3ZjVe2
ZXnj5PHhtECz745cD8tbTHSLyKHS1nSN2PZKvsgWx6aLJghOlfhIXE7kY8mdyZpiB8VLyauFK7W7
YDrmlFaHyn3jUrqqwU4AX3tQA7P9mnHdGFBa+WsXfmQRZhMfsOG4fTPdFQWYDftPvU1+uk9TRkAM
OHbQKPD39GSDWHrX7bWLQ4mkHEVI4B+ySODWgnM5hsGcLrfMu3/FVAq8Wb1TRVqbPRcyFkENXjE3
MWesma2VkO6iyJRAeZgkWsmXcZvU3JphpVIf7WkkkxuOln1R6Jxgkl4RrBbnsFPM18F7SaOAba+b
x63hF5z244KN8d7qupmct547XRFQb25FOVLz64PRq1j6hQl/Cih3/eAccp72p0T9D0/eJBX2qrpD
sFxpIgeN224cArFq8s4wi0i3CnCYXIlJE5j4GakSt3s5WLHbSVJjwkxM22BAn8ah4IERw26TS4iD
D8I0xHY56CRhIEgi8OADqj22h4cxIbs71NWZ6+KtViIH04cq+PQbcRyaml5xQLXHwxcSrYs22KnV
0o5dqHIzygVhlGrzs57aa4991TIdT0mvlq5NrqQgL8r+34/d9VoSgfhUoK0ep05WIgJ0pEuDiYBE
qG9/RsU6ti6MRgFCm+hSKRewaaWj/VUQndLL3+MWaGTZBVDi1QfB+v2VCnZnQ/JpdeFoI9gRBz3/
XajdrNju/wQ29cE+EzPVcdBHSWv7VwSrJmQe5Bwe1P8iohqHD/NP3i67zOKPGnwpTkFgYeUiy8DA
UKIgr8ya1SUeEiil4LSkGYMeqb++3Efzf4R2u3BVIiOaLuC2hcCVVy1vqZtgrbGwvgPdn69LL7QI
EnHUGy+62DW2qDNzre47g+gd2DzajSjrfWoN2qH776wMCMwnAZct9eOeaXHeB+2iks3AdWCq8epP
2ydNrc9mLL+IAnxMDRFIvjBsgNJNwPaA8vck26kJ9IwJCHe9nwlGGprUAeYfSmmcqml8bSEGPWUs
vSTsgpcOSJOyrp8sqiYelr1MqwDJ6DSpssmEZH3Lbqpe7LQBAhCLEDdfsR3CApZ2at5+G+shbCIu
SrhzbHBBjxt+DALOcB8HOUM7Vx2SigPjlw4elEbUoy4DWZ/Eu5dfwUWwLzY5er/dAYnb+dxv/v2X
e97axNPi/GD3Shq8DC7mlbzQJmEdNmF+eiXuFLpdvdm/pp1LKcqmzwhu39q7xOXzAu9uYhsW+hHG
28XiVDOrBaeOunHOQ79xFkDu2pJ96c00bZ+FFgOfu2kB/1RY+lW/VmDLHciTckWtG9mXX5SlkMMB
CtiWlOGbB77dRLjSfoWBpohWRyR/JYoZ+ykqk/+R3qDkLYXsGIwvVtQSxBpue7WGqC0cQJKMzNa0
4p/rcpG3Ck4aw3f79Q7qW2/F/3JF0tpcrpvqhcsRk/YnQjbBsPYvPnh6hK5PjoRNo9V3lxg2ho0p
bJXKTwGzUIkFjW9prRsAcWx6vjiulSKVENG6KcY39PP7riItMXlDebOjoLiHq7Xa9mdBhQEs33dt
d/DttV0WV10Moi6t8gW1W9g13951b7barKwhXLPlBFnHkMUAJ40dOOPDvgBPNVRC6A8+sgieRHv7
GhaLBPC9qQ1dDdrOaHx8r2YXyY97p+Lon32v/yxwA9tJrPFEfGpp44kqe0JQUvsd+VfpW30orXkV
N9nMZXyIygjCOkilt/4PfByFiHNbcxVejcB8Y+Vc4qf9Qt/N69uA93U2pPq6+EajRi+II23FbKXI
ucY1ud7YJrJ8L2ypnwLZqr8oFdW2zxtTuAXwaBvFSGYCbyD77r9Qkis2W096qSkKDKYsSalY6oB9
AvwVtGNGpTpvnywDhw1Qu7G0TzenbIU0pWutJBZl71gd0cWnxFhAr1ipPaubqsVgiR3yedX+E9bD
w4oTpTH8Y2ahO2fwVbUWXFNmO5GNSSHIlNojPvjjrHoMDbYhsqdTYR5ZytFADJemPtTPUz24fTJs
cL/lY/RYYUDV8H0FcJ64tSra9l1odl0L3OBVNw+GOY0lnASgisdcxG+oLLHkj5ayPDNPRUfCAki+
atbd+hVE8E7jgbuJhCfKAyvgfNOP+rrh8Aue2QxpT9mzAxcwy8x0bMzxB3N7KpOwypv/cjxbgOLe
Mp6OY3jppwB6xAsc3PaYcAPCG7asPxo7p178GiWP7Djn6CO8/HqFbxEWC9a/FIPwlDBKQdpaTfF3
vZgi7J2weArZYJh6lM6BcdItIyHb2dU5yZwKBKx7vkr11rccCf8LNLw+kxPMZpVgUfHik9Zrvr+w
qWXYoiHu8LxhgdmtzBmeh0XdKCDhU5NSlnZWXovLufsi/hdTLlwtk3Of+IPpT1OHVS0NF9mtfkWm
dCNd/w0EI9huf9TdvZtfJE/AQ6JYQN4ARdGXwCX31KJlpXNUPRDAZsIv0uidL/5uFUT+JVTESqQp
xRvWQRTgislSrvw8hvo+qFwfQtEHxCO3xG4YGmHY6JkgYWHmoRre43LtA6dIOe7JJPie3CT5lG6I
TkRn3kJHFA/AC1FOGmbzK41xPwJ/TAmF8Egx+YMJVAobNokdwp9P0qmngSLRg2Ql2wataUNF0LxC
BFJT6LKcXrvg8Pkv+VlGlcFknpFbaDVTdz9sChv1QjnYurQCxlKf6L07J/uwKiifBxoTwSo3lu7Z
shgpDCxPlBoTpnj0cKDR+QOp86pWdWiovTw16vJgkuqKRUawoeX0OaCGszwDsB2g13RIGslDlKe+
Lc4u2P97uoPguMmzrMo1i44WD2GNx91CYz6Ajlr2FAIL/Ca47a8jzNrs0ADdKPU4Q0sZaNfYTPqf
A+tF+SIY+yxPvvEvDAoa+udomWQBpb+jfddUk3SoTnMvq6/RxYY1uJhaawvr2rCtK9eCQJPhhyit
i82knpyzB54EHuGYqyLrkosVFCyq9JhOuy1ikWnOL4fW1fpKAZa5pF1Np7AiJazf7k/Iykr+4VFn
t6/TpTnK8B2nHcjwBi924Ipru/1rceIVFei1NLkzyerVqQUG8sCSqfZzkf5tljhay/5faHnWtwnR
UKtvWUhM0koBflE+RX9wExRO4ILmgu3CEydUDNO4KrYC4hatxaG93gBxfc/j4BBmxG3/a7RhtMYh
n9PFyaqsW2zSuOKTMMRBO/dzS2pgeE2CWy3Fg1jjsHVxlOjck08rdI6VjupuzRnzL//v9b3Ebzwe
4ID3FlC7A+mcnmaynhmR6zBN2PEkjulokw+2eg9MHUKwMVo+cvM03HBEA7Xw++09Dv80AzXN5SUE
RBPPNL4WzZt1Fzp13DXpx+vv4+uZjrxJOsmpfdhEERqvIbKOChV2plmsIIQsBgzFNJJxvhtot1yV
wq70rqei39YtUqaDARMbCjbq4/BLzicw03AYeTxto9DZbH3dZd/2HQe2BrNnRVfdkGXuWTTovORn
4M55tzc8G406Yp7Fzj36r3izBXMwbxx1NIdXhdF/EHRqqAzup3ZC9xdeiDAmqUbfNDeEGQbIc7Tc
DhJ4lidDKiw3HBhRGtHp891GZJe2nMhHNZQRckt++gsxKi7pjtHkVybxE1XFwq2K1vLsVy4JNXl3
7ks6De+q2/diVgwPoqyCxDue62mcYJtqftzUgtJXEFUK6h8Dis9sZvnu61KmkpVpURXE4Vn0Yu8C
TI2s7A9nsxbDkF7Ngpo1F0p3GB3ORAlZACT12wqry/sJghICF13NUC/fqvUXmPUOv/q/GqX4N2D4
6wTaIlPq3bMC+rEA0zSPa8hVDGSD0EB9RONkdopvew6G+l0uPsjgdG42az1TEt4N9Xxno3b+l2Kf
WELs4j4MuN0aOpsEyYC+XeqLYCMB8K/eQS2Di0n7b9ZyjA0NwQ9uZXQ5NOv7z+Z6o9H46bDJRquH
0amhQmgb0Nqxu9VQIYAhv9jNkPnVQf7IQKsRcpYpCEb04HoWvX6B+4NQvMa1JCtbDsWutbrHlret
PRQO12OPV7eL2Hqm+V8KX6JS5SQ5CFtUlONppAyv9X38JN9IIJ5Zni6djDK30GptdjP9pTwHf0nv
0C951Ivca+rZSUXpvfvBOd/RCHzsXYEdi5KJg77XAwrXn0rwFBqkQkWEAvqoGM+mKi2iiJ7q3q/J
Z07XyR/wqCbCAohi7M3EPbhGu7nhmcq41dauudCwpZn/t/acf5DrzebXPX4qFTCMj/8tZ8rC5vDH
Me5Mt7JJXLkXgH3QBqr5lKKszaGIYXurcds/gdUEXnVJxzuANiIW8hoBpevEOXu33lpUjEQc2pwR
lWkZ9fRMK8y3yvHzOO0pCeS266fLSYtTTtnQVkLOwy4ftEGCwOGHAkvhPUBJWcepF/pjD2bsaGg8
TVBa8VMjvFTkxxkUr+W/jGZdep3XzdhMkTsh7TRKI7qOE2sdG31DKUdrd821qaE8xHSqdGa2b5c2
jh1aa2QI7UEYyWwizP6agBCo8Vc1a/VEVSFzBSRVDwHPCWZDf9JUtCOeNnEM8+Nwxhx4En1p6ZUq
6jT+P/sbp/3m+qn4+SdFMVdvzkT1xQi21nbQzb8neIPt1GQ8yIHSUeV4uMIU+oehKO488z+UG9pk
Db3lDoh6V+NFevXjr3n3KyJEgrRs7Vt5KX6RON/8dD3hxvobA/KJegwHKf+D12FPruny6YjPm1+H
jOQnqwacsE/qA03bdLf91fe4RsRrJrNFB6BpUchZomW3NemfKlu87xRWdrX7K50uJ4Np9JsGJHKU
LSm6r6QtPF2bcOpFd8cPNt31GVEJwtpzn3uTUC7dih140EwfkJVAWpwdoafamtvPlSAA+9kq2Rbo
uRBYhU3xZ9DBL09hfZg9YEXGoy2VSv0xBF6sTkVJGuOwDhf/siEz1uBIxjMgOl36Cvy2EA5HIGSZ
woPEDY2QGs/I3d+1MAQfRlOpTvsbb83Mwo7PnuuY1lNf+gpYyN8dXX/rMswz9LGzN+yKleRIMQBI
2wVtGHshgEv61nrbd1PSlf962zcU8IzvN685Kumqpi9UTtpk5TmB3rAnp4w8WNxABizzuq9r5yYd
R7iIlaSOaFBqzAY2vApT34BrDAnT5obbvSoqJGT6s9yB2u89pn7eq94zEXP7ckbdHQ46417QxlKn
NyvUwkK9zdf3EmEhxzKiJ2UV3vZX+9IWYztl9UkOJ1zC44zEnNYqs6HBCppgDAnpVkWwb9J6q5vb
wUBZhRG1GrvSGquJhlgN33E3c4OCrOaqfgAaP9Zv1X4iqQQ0x8jevfHGtwVKOGlZ8bP9F2UiYcCs
0XcLOnvotC7Jkme6nzPtFxqSmnBcpanNLj+IMsfToJeHeH+JaEqSpNzvDzPduiF8JsK133SVACVG
qirYcuhebonbkB7nHnOK736tktvOQ4TTn22mPpakfnp8/A8Q77nA+/DN03B9XEKV/ktktTcm2Hmz
RyBIrCTZZuBTnt7BfitkQkbJMz45D56PSOuNHkWG33OESD39U+LYjvUQ6X1lRwajx/2YZuj5Wpdd
Mn5QW/m6yr60X+16bz8i9iOKb+wDGGs7mlUNGIJQuH8MqcMzyzDz8QAh4KZF7peRfqRmAuGNd9Wa
purQ1+ZGQb/re6yscas59biOBLGp4NeP0XKlFWU9P7PHIyTi77bww/ELDjFYlPeph/fvwKz3eDXF
FkVN76zm+tUaoUoiOkGECZi5ZfkL6I/sHIgCrBXHSuY1sKIwRH+FbqlrBZwcB8lhMBr0zhNrtUgb
rEFTOnM7WgX/2IylN+fqqQ4baZNkYQ3cNazzXtn9hj7jZT3OOpM9v71ZAACRIxDdPVG1kHH2Ls1n
xNs9KDbyV6vw4Tfsln/WYxXNZuHFGIZkZBkMEDwVmE6NZWX5uoG9cFMOnBcol2EJ8lGnJVTgFr+S
6f4dodZLOIywHEoccB8t1ymgEpBfRFuDQprkY3cS1uhC5WX5uQYptA/MM9QJdHlWH9rYEFA2rvA7
0VBX+edEGdbvYcrtWCTJpYOdNW2850ydpnadwmFV/oCvrlBCaYoUoVmB5GXKmwfBu28FWswrVGW6
26vq7uhVpphkTi6A/xPG2065WKikqszW244OWmT4bQAnbmBRULQ/VgdBXguwqcJ0OzKkTI2VlYjj
+TdJpVtLBz15j7gmx2krkcvpNGv5Fd7ArPdeQMvkqERctP8ji94d1tho4NMCiktiYBLux2OnZAen
HpQjj0vLGfXoxviysgwG7LZYGqhhMTH0HWFQBpEb31W61tr3skkREeBjfj7s9+AFWI5J/oOnPTNo
QEdfQ+THd32O92J945EL3dHtuuFb0H+vPS1qX/Hi6aZ1iJZLbV7oo67RBGFXa4ldEhNQHnknGZ4E
PdKjUiX2XrBxx3oTuqCs1qBLf9QQpf458pJOiugJKPKOxMG7YuGAU1fLr4lWbn7gUsguySXXBgyH
+6M6gkpfFkrwJCvyn0eN6pMP0c6Nelyal2RLkJ1/gdWkfEL+b84IQ09ybVfC/c5XB12KbBFNBVIQ
EIcc0WGZ/Oc5esJJ7ZGlw/njqJzd8lYxp2xxdcj4pfsgvebz9ygiMd7zVstoF0dEe2rgun/IWkE6
ce11MTAdawI/ICH6xfDs5jtd+BSzX9uH/NYe17zXInNcULOyf66rtTE/iWgz6wgODmabp9iNynix
1j+kR4zRGISnX8Rjjp0psVXkXSqgkapC7tQnl2guUyS2mE+FcWNznbgoKcC+oXmincnQAZMFKwvL
tIla8Z+b6e1uqPxLnLtZzId70aU4M93ntZhv82iL2EimHlzUG3xaorOU4wdSN1iiz3AI/LAm9G/o
IG/SxMMXhhHH48jr3iKexVLlrr4b2mjOj07Uy4ilRWXMUyZJU5Jp0UXMMhx0Ft/s4x4MaUA7Styj
+UpeNdNElxlLJufC87OVOLUZZtqIwGVHztkQ3l0MM8yeadIJG2zndsgaEnHX2OorVqpxB9MugSvs
eO51HVTJa97OhFmzT1bk1A/TYPSTyxL9ciAS2ekJQ8QXAHNFXVoeRJVaucNbOhrkO1O7AsheUCom
5bs64cyXK6wdyljuHZ6oYMZ/d04E3TVxprdc+dvrdJ3+awi2bmorWsG4TTdvKw+n/ccMRxzbkZQH
bcxUTq1MPKWRgI6jhCBtIIxoErJDO7OfqBfm5kzKRTXZjWDjW0uxcqfAqtfVFRB+CNF+hNtSd2WW
96SHeiCGMv4U+V3SQQD9swYrGMWWSBgIKZodkS35H5LrgOceg//YkMCGCeHSGM5QiSMO6Twam1h8
V3HhTdOqNj/7F6eLjH3NtyT/ZPU/by2ZRWWj5YtIU5ARefPMOd2o93g4E86WTI0MDQ+m8Q7FXDmj
ZxHvOyxcKc1cNrn6jOF8pQGciqTLadpzR47agLthUt0kew+3kgo9xhcNcPY3//fIpT8xCKbe0tFS
DF1mQv9FElQRWowZHNgYTXbv986YVgoEOx+eKXifUMNclvAbOcAHOOkoKi5yDtG4UDJAgLF5hjnG
mKJ96bpDKRn2wPA7depyx/d8UX6+nZWGMHnx/RK6dw2j/jyxUlzCiugD9s1Qj2ipqWKlug6f1uMu
hdBB27A8mKHUPKsBw3oXbwKNfWckF5g/74oc54OeJ3xP4Q4Eu4VySHawpaIFEhjaT0wU4Hwqr/r1
6v3pQo7KCKTYORKlVA7v7l+O4cICOCjtDb+a4e+HTI812wI1OJpVYbm+F7/4CrUTrw9RgesKUgOl
W+vtZK+OLJk5iXiBjx9oKBx4qWZDMvO/XSKbCFAclXhpztWJBKbZK8GaNOhLgxr+IFvREgOUNXbD
xrnFM5qAgoLYToZxWJOWQnSxH8DQqYSZk0K2k50K33Rmln9qPBMqhs1HI+yDi5RpwAJgwnpr1NQ6
mP4NuWpp1LOBAZ5bIxAH0JfCNDmo8rFcJ030G2yrjDn7Ysk0MKmmoknS1QLELzJW7vDT19O3BEX7
V8ozll/lT8Zjk8VdfkOwG3m1NakLUhLF5JcRbC4KmaDy0bmCeM/QZijfDiUsKb1S2y3ND/xhX/uI
2jsRKlK+OKKfSQJMrxg7Lnk6PebA6qmMLnkZk1HwpHtDEKYaVi6JPjXGrUz488qfV54Gh2TG191V
bvfiKk05noRltf4Nd+Rfh8ahKvGmWKeIcUMFvAVq5+RLy7GJ1SzvyNnHmQa2BRlW4W82pLAUCP+s
N+RvcEfxiImSEA4cS/iBFv2DYCoCoxhlRVQ+FbOm71IjmTeCYi4fN+tBsXbV17JuEnH1rJ+u8fZT
FYATFnCm9dnG8wsBVh3zgHod+ubBbX7VmjpPqjrHHwJuKk4f6GQNQMtbiz19BQXuREtGAlips63b
4ahTUXHc4bEDCYQDSD/aXKzUzXMlyXRZO0rR+5bKY3yVCWK4IQh6sY70rm7kimbXN80+8d+EyN6j
nycbQqae/OI6cGSt25HOHusdKY3GYNl/dKIeafS2DkH1B3AknEHb4zTtDbvzEgfBZHhJ6olAN5dp
Nq5GEq6Fel+oMUpZWsYo8U9oAJfJLEQBg5tgE7Nz/xJMo4P8Gy01WMe2rTdgqRFqxwL8usc2EYg3
m1f616IcUNDlyCQkzPoAUXIo8JeiK7sx2rJWPKEk5AnGygL4DHnHfTPGsZMc/WRwkDWhKEyQfsbV
/oFcDjMRWNmD3wPt61In53pVmx6ztbNzNCGcFbSbXgwEWDNjjGESYgr+7nQfhshjd8VpnsiW6W1B
QoyR6vmO3FuPW3qgynajLwlNOcj1UCEhyvRbwtuwQIT90Mv95rjEPFr7cQpBagjxRMxth2bB6X8D
xtsJgiPfWiKT90PWldi7FB77/3WF4ixJ0X8OkH35BCDuDuOO0ijig1kfNjwx/Xz/wweHk8zY1ZMA
3kF6CZP1J7YFby7nKeObmJbQIQ4uq5pbKI3pfreGlj4idI7iJjA2fbxiU4ZlTCDh/fmsUnGueZze
M/5+JY0MatJTr5m41KS2SWgf/0nS9jcVtePpmRg+mLETNS9SnwYNrLgiWD8TqEmE57/qHbPFuoDH
NVfYsITcjTWzVoNkgs5FKvo+h//1EHE1O/P6Wif6o4NeI4N6ZI94urdoyWJ0AmKnJKI4vRFyq5kz
NkCJRJbpA97qwGzXQQ6myrTFzAG9JsRiK5vscTdVvIvJ0XXez6503Cvlq7b69ZmNg9gedyjUEfD/
BwchBWj2ckDCPrCORaHy0W7cjMNdBSQ0e5NB1qkENzZNoN52aIL2A4YK1dA05hgzYdjkg2YU2Zv4
e9t++vFrIXBdc3PJDx41ZkUIBX0bAhGAqTOnkrsSahg7kLvxyOP7VpA5+UiCGXf7kHfuAjHVFoks
qTvR3heemkEWVS2IzrFM2WLc8CYhufdJgumE4OSyEARlJtF/VEp229ap98x/YIeI2PfmOCylRpw4
66EOH4ZP3RT7oNfPbSAXagfE49oyZkbTJXxtf4huZauBnfLtu4mhTgCkGjy6dTGYIA/B5vcCqHDy
hx+5kA3vCFsGLQbswj/FZEPYFqOIoGCTcwVsAWlvLZiGl5+so22yS5sIQhWzGY1yz1J/era8a+sG
XiE35LaDf/rxAs+xaVae+tvOPFxQUlaG092jdsYc0jjEbY28q/hJ5mKbLGfhKtmsIAdNaV54YtoL
dVJmQ2VzVs6Tes6u+7e9h5MfHZLt5/bC55l/KtWHNZDTvLu/LzCJabODyml7RG4ep44etPv0BJzO
CCmOw2R81HjBBfC7vXDbuvu/iQJwMN/tErkmF5kqAlk0Jlw1T8/nqiEkmU6dy+9gVKs6e8ybqJMZ
mtsnDFSWe6dpvRrQfkh2QpxWS1PJZ2KX1aiHnTsMXkGrwuXN4ka5r70UgvWbaDCvR2xcQ4f7n4aF
nmAhtx1CvKLNssY0WvBsUlZnajtG7wLoNeY8GEOZ1SAQmYJI1wcqdTVgtMWVnWh/tLIoJXZFrmJw
ig3vl0eT2QclmwCZHXjmydDCO4vYXvO2LXNL03S9G2glqRdyIW4dCYPv5AFKgFp5gt+yfqkgcxpo
q9AhJB7uFRWUdZ6IwVrFwlWoNQ0E9VnvPN80+MNzLncdxe1PQrfnr3rNpZdTdR0v05FctCktmXSm
6OMPg+ELdXjdBeeuCdf24sglSYJYlWMK/RmePg4i4b+kGaMvJ6Jjt2aX3IbTsqgCPg5vtF0TVHP5
KNs5vHd1KKzV6drN4vxv9kTDyn4986wfSnBTU5jzCj85UK5gGBSOaOOdfdCbAkT5k2b5t08s+6Ri
ui3dOz+uxc7YPahtiDxoSUqRYbvT88fHc2SXnJmxwX+bPCzaXagme4NwCRL+MQVjvZ0z1qwJOUt8
nFQsQtZSCuzzXjBhERrwva07C/e9khKi8ojq2QwxETKHj6TviVtd+y/Gs5gU1KRd11392eoMkVs4
kOKGVIHB68K1ecSMTNRhWo6tE5to+rTRn4fYfSiJvxGzancR9hJ+PYhb2l4z/WXsC/OwS73vQtS0
9d9sdIhbHh+li/BjOwo0KXqXSrZ0SKnE1ZPhgALq3MkwWPcWvq2QWRM4KFHcV54HAf+hCDE/HMrk
VaI6wlXQvy3pyhypCcp5iJ1l01HmAq18y/To39ep3cm1/Y4pyYeeQRE8n359dR6vEdJFbm0pv4Ni
Xth4jioxm3NSCOaGGd1C3piSP1BW/eU6ao+6VGKfuJhY61WRKZgFe7CDxq2awyPZBKYNy2vTwPpr
nsZkbLzakgCPB+9451UUMHxlllWQ0J78+Pd7aMnS+py9H/GxO469arz/HRAV0I5aDNWZJ0JBNftr
TbDAW5KSwAbUV1Z997sy2QMsILUpnP/aUxKCpqrpoRhgALO7NNalRvsXAnlIsCYULA8Cnz/2xcsd
LGKVKF2Tf5TJQZa62/bEpBS8zTYbPQYgHPq4xZdUnWtAL+oUvL4hoSV1/Mj3/y6iJvXB9eN45fHA
no/evWS5XAeEeClctz7AJIJeDD3lK2k+0+f+x3rJQEWGDnKRRmwCmMzTzKNzVbgzKWww/Tk4ln+n
L7uQp98gTsVW74tmTs8ngb0wADi3hPxN0SiaeopmM5ci0aZeSqyuN/Wu5ccHTLhIFn4QWqLqDJIE
dVElAg7XPpBRQ9RzlwgolZ/bDDBT3NpojXpi/mbC9+oKVAKjqoMhbjib2zQso6fFzGCpkluU+Yjo
5JKZjoCRkJgtkY8D/AkwiGCZ7PYfRZnUHIQfjfYpV00VOC229BvbxVIJUx1If9U2+caIhrjiZek7
KNLq6RkUAIgAqWG7FEc8hLT8D2jBww7bPF/0LMYwo/Wtlj2Q/OZVZvKVfl6el84P/NzY0Sv0ug8D
1yAvTBPNOm1OAUBN40T+WqFUsATc9X4QsPvQv+tLf6+W1ofpIzU207hWKgowDFv3GVCQqBy9rp1Y
Sd25286ocntlE/FEMQPUY7ktIgc/v8TmIAdZzy9ul17wAI2NlFij6RRj2KK+dsDjZpbmOdW1uSEz
Y4qa/hiwFC9N4SAoH0n1CblR0xli202Aj+ZgICrAIqibEwfnqkM4MhCnygfhrWsG2iFJTO/y80in
DaoBI7Cag0hlIyftctUPyyjvHycopyNKYgCgvybSOuDy7xkXXsOMi+lKhjJ3Rp24Yd72zKpDxA2h
PVPbhBDFv917upD4b1ecM4lrfdY787S7XJ8yXlEyTork8QcTgDQ6dgLNH4nILYVctT3fEbxikzqF
P0vab/n/owNka1kNbRQ2LlEY89EDQFvBPGGkBySeRYY1IA816q9kws7EUhnz66weo49A0CL1hcwg
7qK+y6j+HzxQELCvrFrj5s3dNDer/xSOb1QbOzQ913tlt3nDjiveNb56Ur+GZqPNZ259UfouDqR+
H103xVkXf+rmrvA05b/5qwiaVSMWvp/u2VfVTnwzBhVnCB0sXhTqy3yEJy0BnrgjC2NB4bzdCXdt
ReoHkdV4n43XfNyFcfgadeO/fg4KDKn/nuFwOLnjZwXRpaIR9GCvO1HpWAqNpMBm1sOpi9L+XAn9
VP+Y8S31q+i4QY1RdfEAYZ/DufhfTZud3KzNloIxTNayg4Cnj6+8S3PsKaNgqJj4CiToKUo58fNH
T1zwHEk7lpDJBpCZ/aaPLRatv82zfxk5Fw0MBnJEUuGfwe+orUmAGDC0zEoV9jqsviGvhd+XzWue
uhQHVdkwjGjMmSIwiq/87g/QVZDBMV4mXfcbUlaVDCogwzbDGkMJQogoH4lhjteQd0qGbJd4rHz4
h3Hqdtt5+Fd9Yozz2iElHOzgcbEN4t2+KcdB92JknXFQMIutiSnMLz2PMMGkPQM5DmnhkkeDQN0X
rYtUE1oO1Deq/gkKXJAa3GGaLQZWPXnieUh2sxBGNG5VUconMuaXHamX2fB1endvizQtXd7hNQFt
e7hWdI0OLnuvOMg9OzQv5sg4aSHWAH8mLEvAS9WEjm8jg3S/QTku22HT8+NYrZJsrCCbbTF2EOUz
Mm+jZH7CYuovOeO/HjZ1AGu62OU01HEHwGZqRVau5zSLgf+2+YJftE9ncaq4OTF8NrmM20e0s9GV
QLN+aSy1Ak5cd71LZrKdQilZ/neAuJI8RL1H7mMkGUlYL6TPoTzGOWQ18Qs0XSk5w6f2zsF/4SQ/
ARKiNSY0lFh/pH99twBh7Aa7Kex0seAeFOKmA704rkkJYd6zxVomuxOA80EyIX/2ts1oGW36JoBa
PAI46JYbXU2j5mqZzW7ZEaYcOwAnh/1rlAhFyF4ZwDFKE/hTo0/D1bxiNzdQPDHDBoo3/4STRykU
m5W6UH94oWpNc1XLIgtfA7anjQ6u17CGRQJAa3Xkk7OIuPg3M6IAR6Od+KxeSV1zyPsQqw0SASNf
XrB2I3Gjp+1SZZsoW10eWwdHJ/5uyjkOYsVZaOGKTgkpOvDJ0fa2uefWd9tat4WKWPm/8Xr1ioWs
nWM1x62xqeHsuLG9QyxCSt7vGQjVojJDFb6MzChnGT0xTIjnndZ3FgeFTMNImh6s/1waRiwcT8Mo
yqVq5MQMUuPtnZdnMdtMCSRIGXocc0hrZ+dwR0pHHnLdrknmYuRn7mJJk3y/ZSw0l874rKuuMA80
kix4xIW3Ej67FzvY5nL9owli8xunGta9P0B3C8h+4nz6Wn0SfVeKdTMOapI7QVDYhfb1sQmbnQjV
8RuvgTh6eM/5+lpr925ZhpxAWxWPC5QqafHioVEJ2KXW6WmiUz4uPFKC1x2qgo6gCXn/jUxrTjrP
j0/r1CwULjMmcRF0dlY6trUSX3j8f8Z3cedDP2/UkU6yvVlm0fsSppyGV6xD7KPlmB1FVDZZcHD5
4od0EukQfydchvfzTc8bNlJFOACohGlyvlM8508RdckT/irKrkD8TCKJ5LRvK/R7mJP6LiojYnSH
T6jz6K2glDBD8QKNHmoRQx6QNPjpX9l6zlSpwW0vI2ByaWs6kM+JyQ3+IlXPLA4Kdv23kkls+0/J
YzC5HUOPErl056SLq8xX27bKVntyIlUVqIvmaUixiuSryJ6b9I6sKg/QrYe4Ci409BtZgVtmup/S
ACJxNoIO5RtBNGGTHDj1tkQ/BJZRpqYP8X2fAVRBQMYrdmwrwGQNJQ2EsGhc+B1X7DAgPIGLkALe
DuwcEKdQ8bz9gwgdsD3SbBtUvMEpwQkKQ7ZXFELctqSu9B5meJMd9O0QSDurfIBh6MH0DFbCZujJ
idfRLgUMa8Fxyy/C/nJT19DrR+ftS7dCMoSmiWG7CUz/jOPGRJyX3n08KeiHZh0BLYPIyxvm6Ah8
iGt6P8OmfAZwXjL5jKEu2W/RLZdRPGaJoQXTraJFmiXEoyv+GHC3xKara2SWvCYenIRzuGL2F2Gf
thrRgnwWc1iYqTFSPRUtg8WuRx3HcnaypGf77wMfKu8uMqkBRkilEcOsUnm7zdgsTxLJ1jlgs3t5
gQ2eZM2A/w4WOa2Mrn/sNPFUWVcjS+SmqGFHiR4RtiQPs6ibqIX0jg+2we1YIogYf6876Qa1VNfT
DOF5MdKZe6+96CPJilvakNW0DGPztg+mLj+XAjgLMMFVjf5NMjDMBQsl6zl4yTppa9qExfPFry6X
Ol/I2w4nQtjkJQtWdM92aGxdf+VuS3pj3iXdEv7bnvps8WXiOU2F/EuOkF0vdjFymbDALN7rRLRk
/RPrFV5J6NIQM5fyUBAIcmdPmPV2s2vZ0RUrGS8zCezUwuwiaZb4Gs/UUSGSCTZudnX3+oo04hQR
ewr1kTDmvUZWFpYra5ATmEYrOA+FmolkeYcU5VLcyvSwa23z86q+77HYSrmTSdWrpM9qkh+4MB0i
hvHqr3JOqLOEamyAVvx0xKCIA3CvbJGrluZStHN9X9chYeKKsi5kycZQ+RL5YKm0B4YbwQ7DyIEU
EWbGIYi0hMlDuv1QUtWbAK4s3Px85IYoVDjyDlD8PJr/WE7LkrvQgc/WKpX65kg9RTINQfOUXc9Z
xDYy8j5FOwJSr83aQdl1rrmSs6npL3C6OP71t1QKjjqjf6AfWywqlbZBwQcXcesYdfllO0y4Ouvs
dJiKOa+r37rwJNoBr9urt0uja6h7HzLMm56H+CDZbCnPBFORPPheYFhgG9miq7+yv+Hns5/fBj10
dLBriwt3LDdSxthQNKcO8Eg7LxFEbN8zTfndXEbhHiOjCITX0U5vFuq1sjW2CDHIZRfFNcm9z1uf
J+4KJxWstelLop/3FtPawJsPbu+MjfeWei18wwsK2briEpl46g1ajeMD5cHCYuKsY6v42zBWHxHO
Wl9HZRhbSlCWS1JJLc+vJOv0eLoI4rwfUKnsyiaiqdo51Tp2Ppx8OlhSxPba47yxi2m2s5rG6v6J
/hcHEH4B9Yzrto4SthLAWTpSv5Xxfmxjaa2f5F3WwIcV7csiONys9rkjGooKWp5XoHk5H7eDXVLb
8SIX09BmyCAVKVDD/g4Z8OUSveEIs2WlOEZ5pgHf4g4UAks1pW4R5EkrrvRUeShnpQbpqi3qwJ7n
9tYSzG1sMIVZs3hUmXZFrYdfyQjZg/2+taZR4GX6TFPxFsPLYwDYRYx34VqfAywiI9VmGcjcyozP
6waa8ROiHnAmVPEvNwLW/wGWfL2C9GHphYcYcWo8dsZc92i/nlVMSbdKey1SO7wV5BoQBbjamLPK
9JhpZwyC3OnW8noB6XW4707RavXv826/dxhQiQ5R1J0sWhkYEAanUmEVn9bTGd9Y5NyiQFdoI149
UGEIVvoDudPsaTlYrlR42sp+jMgRE4zG+7mSPaXWKCfkrhGKQxPljlaQKh6pe7q93wg1clSelxWQ
z5c3egijRqvf3CLKiKVmgKmHySlovxzracccTJyvuDj0faD/oXrt/hSwtzlgE/6JjVR60YxVzoUP
JogNDhD0KKLDwcaQb2SGd/sbP/PaQz2jyRKK39mPaQEVoFnXoFFMTP3MFDCWT11h5IBm7Ly//2V5
64bcuBLTUNcNOs0HeqPSqcDyXVCe/X9GlrrDvFNJMjfkzi3/ymDexD91z2yqPJ/CcWbBc20fErxB
f1Ze5ZTVL+0Oaqd3ew5shu0mwiSGAtc0YVw3jVH8j9+gm8zIZuAbQN3WJ3o/hXSGF6EaBy6NQhQj
sOf0ncNT86+XsJ8lBuFCTarl8dQo8EfThUqzf6vkG2eZtwjwSj+JRcanBqnkriXpvKgFD8PkIklv
+26SB8Rc7Ot9tRrSOeemAnHXMlu//dXl8UQretjcES6o4KcW+ZsEwyKH0GNNgV4bYqodcSbMX6rF
s1Ev/3eljz1O0y3lONz8+8geweXfMjlctpQ6owy2px/Php/BSjz7AVk7bfL5CoZz9SRU+gjNfmxr
266VN/mSqoH3mGBZ0r2+AdKL9In+OsJJkhEWc41Ep5RK+KdjzFyxwX50Lv6oyDFLBhpf9hqc0Ry1
9bWU43r6nJdr3r4uIJmlP2d6g5/LLR61YPI/Io1Zq3WkpaJF7EnZjUkeyBtPvMa4KZw9trRnFm0L
vImFzJwuxf+P01PhDQ4+6wZkAQTtvxJNIJZpEgIQ2w2hhLApYY10ToN5XqHOlJ7vLhc2ykKUjLEu
bvJc+qmj/2JYxcSKZuH+85i6jcdATvHuA/Ga6Ro2JAxaSePjzNOA+B+SwnAKNqBX5H8sOWH31uUD
NsWvxTbEFiZpzEgCwZU+dhfJ/F6UCRizbzRarGOJBx6vrwyRvr+8e3s01ZzOKO/+I19wgV5ff8pz
HzK+6uMPOyV8hvT0GbVbCkj4jUTBikbBTTCT5SNc21+FVsVPHmE786UYAHYF4otS/sK4h7avAnPa
rAFXD1+yiyrQyWSkCzt4grRvsiyFxPpUqaOCRLpi/OwtQ/fXnaWUE1jv/PLs1SQYQQkArQVpbwIS
DB4gyhiVIBADWvEYgC2UqKG8Q15vMQT5FWK9ObOjA1vGbEsBNoNdjsmlV/DoG5CybUy14rXLJEk9
Sc33tgv8Gm3U35F3pbmbIV397ZpECcVZS6jBmueiIP2WDqOFFhv9u9icB8mro6SwjR2BFNwvJzQc
QJ1k7/Xf2VL1jQACZ2mCqAwFbVjtTcszCbm1pfSk9hAGnvUBiWdPAMMfh4BMCiFgqiVzssXNrOa5
WXEGOUqX2ADuN5Q4DNOu20NxzzPRaogIoG7vdQ4rqdEYP0FXnXJfqA0C3uH+BiunQP53g080TWGx
RgM/KPH0YCIhOu+NUG2Sx6zTd29b8yP5f89vl+bKfdsopre5r27yc3/4GQcHpE/QVcOqm+ruE3eA
8kjpQz1HkgAdZ/2C6iIQvCdSNWieozLdENcMAaNP1nz2fSty6rGhe6TznXS0WfLN3EFmztiSudJ8
1YyJUtcUGNPgryiNUZI5FK/oxPgNm90J6+idAxtKKQBBAIoylsnDYSIoBOHg0BZDp5VnRPiMQfPX
Cfr7dSPoLyvWarQLjhV5mBznhE1QRPNikplaQJNi1mRjJNul2AmJbhDEM3P4R2gqNAaXv2cZQj3t
wSMw3bzgCRdfM8F3zl9zxQGujISXfzxIIwsVCo0GlRPfF1X4LplFYZhGfcAKo7q4KpjnwHbWwuUk
8ZKmPmFERmGShmMWBL5ElvxsgA13GOhBNhP7oG9PJX6JkAU6xxpZC97Lb9c0axp7kD7+6O6iyYq8
B85ehAnCJBQb3vIpdGbVssNpy1Tabsl0nbFQDNSdX7oAiavAEaeKASHV9KG/vpbCbd5RmipLhAKp
blIA5bEVtsqYJtQPnLcD79f23E/W41Bl28YKrU/lDYRHCybgqtvQnnNB37zaDkFvuys7npZEVoqV
rltgVXcfKa6wAF6zWVhuk2t7zkJZsxQZ+zGpzJCfGXk34R0VXLvX9JCwdvDvgFURCv+aL9cBm30W
Rd1gJLoRxdBGxF0nvAG2eJxeToDGl4wx+4RTRWa4SKgJK7B9EHkUmf7xv4G5p84Mq+hgi/Z9Okv8
B9dDl0b9pYPFnr+B4Rp+zRA8LrwkwtZSQPRg8fcsbCHlceLoIQYk3GsAYBMQcaqpMDIziYw6FSta
u1cKsCbHgWvyvTadjOR4LDpQ3ORHd+2aVXuT695VRq7s0YFHoQo/MozGIAhBzgSZxIOWnRzPs0zv
poUddcPwQPMQ38uNV48sqrF+DRLmd3ELZo4RMHuB/M00x2XoQyl+X2R5JA7ZczCSL6Lqm+SzzrZz
viFsyFclpzfVglMeifcwo4RA4lEcighQwejzSZgNtV3mmWwt6n/5oWpvkl67La5FKDlwtp+pZofO
HLwoaxCx8eaWOrFcvUkffp465zPXf5/jz4DkyqdyV3uYcJjsfU5rF+Amt43f09ELCnq/ulD9eaJ9
YTL8YPAs/knmx+/WkO0Lf+WU+aVnQ8Jj8zKqGELx9DqfNO434+7yvvjlK+mLJVP7hZY5DUlCmYo2
EUovwtWR80cbF0WOanJl+p2ks+AGJAqcD/tjDcH4mLVVaDWQRMJYbXQwbJXRyv65aAqLbrSpqU2b
u9Ua5LMNQYafOFwEPj6QV4+31oM9UbuuXIHqsLm2QM9FBpIVfWpiLLj9iZmX3b8YxBRmHonG65td
q+BZMqTOZMbhECfCucioRwOw+KT0G7i5jQcyE2HpuDGlHK/WRcS0IxziXPKoHp+tGmvdxbO8M2MJ
p73BrM0LT4dNg697inBHozPmO0hR0Sh3SPUl/WOoJhBck+H2ztme+/nvNHFYhI8SdclnC36qFgSe
TVTD/K08wE+DPaEoCBZZrDfWVggbzkGwT341GKV2r3on1VNuuP8lJxUljDSAKNfms3gROCOUocrf
b8++UlbaWxCWZZJ5z5A6d+dQjp4ay6praqfcZiZ/rdcecgAjCRo9c/caIN8FeToon4S/ufMxXK1p
zjZaaZH8mOfuB9gb0qJ098xWaeQJM8RcytKNkZojgs2Dw92Zdek4dzRn2HENYQHDcXyyyUK6R8HG
f4wJnrxBv8mfJqA0a1I/Su7Ken4BkO+3TKtGnXnXmzBp691wyrsICDcKLds3VFJgFt5RpeG3qykb
M9OBbRKKJSR0SCK5iriodqI6WLJaWnVObV42S0EN4WzDrVIDq/kwwUMCFIZzs07D0oy0fY7yT5yZ
T00I8+R1RhXhDiEXcUAY1wRjtcwzjbATE8I7imSQKP4AHY/HYDdP4FlwIjnkAp4+SN0SqFMOfUbC
qF7feMq7Clt9DowidaiUQkqmekd/rCiGhRh7GK44djAYSJ4u65J965viTXI8Mg1DcWtunXG2vz83
cwVH6WHyj7k8yX3DdSR5Ztdzy82m1qb4sxdWqf9VYOuUnglrSb/DKdxOJ8KiHTiUO6qhDGkv/jUJ
63ZwlMKgD7s7qxzX4CzwLs4QaMw6BTIgC8OugoQCj9RtgZtRkkZuijqWYRGKaDxgXysjRFOD8pVw
6s6PsltkM4rzqVSZVu4aQF5cUMpIKbC0orq7joamgQe+MQ2f0ndCsg/fnZXBStj/UopFukMG/uZ1
UPwEPbFt3r/cpR3gLTsaH1n02Jk+ffiLh78h98hoAqreGpqqymxhcUZKCTV3oH2NhGB0f99LyniQ
s8+aCLBcfm3SDL2i82pS4VwvsanYcDcmyovOMouarmQj6mCorC9m2EMd8aprS069AciVPTJnOAZ3
jwnCO7rvQEvjj85KO8cGVcoX1oMnux/UdUEwITUlfPfO9lkXn+SMnlQnPIZA5fASz3RrCVLpXhDl
WyVwjiYq2cNM5Z9l5rAD/R9lCZFLyyTgLyUK8/Ra/UkVUSGBtmqJZ2SSa9fLb8fg2YjFd7VoV5vb
+Y93N5yB6XlzueHuISV0QaKJTZTJhYNSg0QpEm64EEAyBocZuVc3cUuKXcdBFiXacQcsljvIY/3x
0cNcfBBC2CCFoJQ7NAhC3nAkVcZo7KNW4KUHhVCzbuvuz/bWQRxnfodGBKA2hef8WIF4TN8V+S60
3D95z4wOQHYwSSXu8sLtgUC89/M1zTfvwv1XWql3xm3keuTIAbRplzfNlbvkvowNWwrfQYG8ZzqO
HMUNeAPqVq+drSE2RZxaJv2WIEMt7p4BlAU+dDS1xuUp5frwB0EHjJcazOU3penpPELnm67R1jFd
xa1RiNwqD6XcJZZA+AojV5e+gZUOWf+4iTLzJTLwZw58PboAmzNauqJrmKtktIAHJgcXJSEn9E32
Ha00fCCvIIBFJPIpf/dHtgQneRTNInWPGIZCfcEFx+zEcyp0dkgzhWoFJFnbYqIWMFyXlYpbLJVN
9oSfhBUo7GJZdeLH5dDND400Sa/ygJDj4y30qllFp1YCI2CKJ2JagIDQFfPmI0qcF86KCwY/vr7O
Em9g7Ei4CQJm3IbOL37a5SWEwLFXGa7+JKIOnevRiw8AZkiPdvZoZKv2+0gCIouHpTLUDhu3FuWo
b0T4+dPQB04YhbtdnjrY609AIt6VjuWUc9+7HhY5D8l71TZgtK/+a4cpeK7gfDKnGR+LVHUq8vGC
BkRIU0bBJ4AM9qe6RJ5jqsaHVqTaEQrUUgspUjexY5SJh4F/znhG8BHQn+ztYMFM64kWq8k3t+Al
ArtwwYx580ujZE/di7JAIceIb+6w52abSQPIxYF0C0pwaepF0EXZEwUAmZHVpejLa7sgpiLTl6ro
eckljVOgxu/lBSLuQ/gz/8byKlZch0SYulejnO9z6NAzcWBhpWUvxvBiZr114vVr7//uDnJhBdsO
qeu4LcnMgppwLK9o53Hn4g/utM+1wH7eOyT5hZyzgRcy2akXv2lop07xE1hFGCgo9GwyOvziYcUw
OSGmzGurF1QGg3ozuc5rTEDjjPvDJY8/UCzMuoZvydkE65BnJpEIvBxnNn0QUIEnnS+NguqDXtes
/nwfJikWJyX60Rmakbx/SNetg8qQujBFxPl0nNN4HATyLoXkd+Sz9XSdn/IaCV5ajkY1KFg6lmc/
GgksBn3hoCjtgJMXa63Ct9Y2rsy/GKH41kSjU4sRJw0iEWthiuIvD/TJ6ndqU/jN0Y69ePq3LQMQ
c8/K9fDYmAkXIiRZvg7G9nQEaS+aLaN4NsfVs8Ot8J8q6sQgl+nwc5Hmnc5qjZz1wKsBda7vsUQ8
jrOo3jXofoDE9Lxs38B0lupq3KOA9nAAOZrM4lSNq9lt/+3C6D2+sxP5yrmPIzWTCVgCDrXTn/AC
tsZFJ0TvXbJGTY0v11e7J//rQxcVvhlxYTGF2MayqFxGBROTLI+jaO/ps994qqQx90NNcFajs5Cx
yvoJUB22o2ecyZii5qH0ft6c+gN5lF4lOGsElLXrPdUZDXLQRrqITIN0aQ7xET/7hD7movHF87yL
cg4WoYASyKc3Nh+ShopUG9nsmm6ZF+Uo+mO0X+5vss7NNLEVbOLuT66xrFXqS9sKZKuiou0GW350
W+Y6BNAz64f176bzWQDgvAJSYE7hJdcCTy9SPuHhcCWIQG6NxjanMBJJXKnovRxB3DCvTAq79vBz
3gFMXF++ulFATNYg1wTjJI0aeuczf7c4j80Fx2W3Tlc1yiAHLOD/Fb46/ECkrLMrxGOoLd3se5pM
hkX021hs2cYJM9DhAYsLfWvs/azP6gm4nLDZkCfIifXldN6KbPWx4CZgXS2kUS2n7rxE1MTKyOFL
RxVo3ibt0Vr+uJaXRHfxRYPNGPkDmhIoOSPU9LwWM1mDR9VkuafvjayZ0EIfHZ80v0UTVQbEG7Py
bB548kdMSjyhH+dW/l3CUdcz/tTn2d2FeM0JenAsgARXLWlNtUKZQUg1pcmXuyysAUc0oT/F3UGu
xO3xzxpXeZIjOdT74YXeD94T2aRdwXnziM9zCWvmnV4ogXqVMDuY5GkS5gzEPPhNqGWYjunIQX4n
d2xLVoPBPfKBPwcEyGWukdXhKO4BffGoGAvE8ql6pjA+kAoTUNulcZG3Ua2kmNJ7aKRX5D59YALA
B5cXh0NK0UqklVeENA2v5wmL3QPa+4eqLStjtnJ+YQeL6jm/8dAYzsi6/qlKdskjdwE95akUz4wY
2Io5ib6T/2WBoMLBlbzdVUtiioXc2heeqPphV8T5oJ81AcIuFIlIwirqqsYTIwQWNMpY+1NDFWOp
Ae+x/aqiyKv6xcK8QdmUIYpfNGNM7CWj6cT9o7mXh5KvNOsDZI2dBBBcFRZ5ma5EcvGzxvSRCkzP
IoRKNLHF8LVMGVJyRa55hM25scHD/LXIg1GkaDuZ1wae2dQ1566pjhdKAPqJCOBk2aixGjsNM0OI
83qnCLPoJlRftrlqqh7KXyZACJfZZLc5024x1hgwofybFiGhWTJVIpKnDIHhWWqP9BocE/gIm5Sg
QvQuqsONFVsgykgHuJmoAoNT2Hi1XTDQJ2BhNVmbrD3AiBRVjB6PyVISdETX2jRfk2eHOrVlJ3Iw
0rLRLR6O0Bx33blELn8HIHJCrrGarun+KN23fIv/rWSGeoSW2GoKimap/l1K4lmgNUx71INQP1Fb
ya3/qBQYAkk0xdaVNOk8t7x3R+16+CwwuLT4Wgt6k/cjSh96GiIRh8BKYvBeF9AV+7IalSuRBKUG
ITjQcpygWHDfL7p3r7j/WhaxGouDA9z636hPEZhM44UNeWXm9RNWulEze0JrfXsIMKN2IEx3AApQ
JiIpmgGRL8bAMxY3db6wv6bX35D8hqk5R1FeHINzd3++PPx5ibdJb8m0TqIKraS6L4hXQTEbohfl
AUZ8aajuDM1QPxgyAnftdIm9pHtnQ9OQ4+c4AzGPt4J6uKymmpFE8uKKVcrkXI8634ql+HiEI7Qi
o4UiVBAHQ1zwhLQBsoxCQh+/LCbAaJ+7anEOaAsmQdDPCzEFZWf5VhP0BfYLA0QVnX0Pl6BW1GDE
RjcdQ94HnkTiV1gwu3/XRfD0BYU+Z3iBw61ML52/T9olQTC2Z4nE1G1rSGI6umYpAXbq287EmIrn
J2fQXta7O3JQkmzRONxevhmEKoP8U/TeGZlHxEgGgSQ6bCzMCn7DAsUvtlnSRmNkT5e/V8fwy3JM
n3zEAMPYmKknh53uFwZVDQ7w9sluvOiRLRhh1qxAV1CHywMe6WJG2Fl46g5NT3vwnHpuFJI7Ilvd
kJCRC0iP/Nw3x2XY9w3BwCmKCvA3SyZ9Ljxjee+bTWTPSRnbbEf5JjY8oM36DVKnGNrtc30A3tRA
Ksl63pPSTibm50GnpkR0g4VLLEsFb0N2mPTUCPFDfSK0tAf19dYC0gWWV4hk682SjQfwtXLXKQqM
NtUE/ZLXNvQLWatCvXyh8NG+KvCf2ywggIpEwABwKtGMoavm37dgjkRkFP7QmZMuDNz7SIsiCKJ4
pp1qOuzxpPs6qkcoHXCVcenR5fBjejiw74wGfABOhEqapUPpPbquJRW0u0nw2wps1OdRHmwzd6xd
vEnKsfqqdfNyY1YJ/7UWYC9o43fSUZiYLJz/+RQn/SI3V/GuDLLIuvUrqZST2x5MZUdSLuT09h6Q
WCqhRy4KEjETIVkh7SGiyWATR6qjpRBZOsbTpeXo5OXfRXmGlaYgniLP3XRFAUdg6PTsDnwMnrLx
7n1WyjRUFJWyBKUNWOd2cT3UM2bAxXUdCN24+35V9QqpGhwtsKSOCCZUtTXgfpex6YD0NpwSUojQ
lVaKQFuTYYDvdEArFT9qVS7rlDQKFUrj9a0G7HF+z3WsXUDgrel/GKEQkZVe6vqG6uOys1+/qvAs
QywoAF9AFkKGscEKwIN7AghTbMdicSX0+LkceM7dvZuSCJgFfv+s1MvrlMmdNAPJ9hWOmRSIarFY
MaJmo5DbuQzE3A+R8EgantfXZH3GG5B3rLyimKR972dK84EmBKqF54Sa4A+RyS/qoBKObXA5i+vq
PMTZJkHM0nHJVhe/wEvzbhkPCQr3fo14mLsKUaztvIZW/jwQXNYbi3Jh5hzKHZx4OvCco2X4HLZo
ek+ZaLhR5S2eqJr1xJ85M5mP98WHjevM7t8ln000VLYj5VJxvkWPpZrMcmHL8EPLoLAfeovxvWOM
LvT/iE7cW1Wnc8djA90OTVBbe8WSDEVbGZDZcfakrqv+n1R68vvStA9hakAGKdUyxt+VZU2yxI73
RUzxEstwHvAruJ+nj0zH1O/TrIy2b8YAKC3JZ6LhhKq7ZC2bV6ORJnJVUJtF/9JrwIbMJTleILM0
k9w1t/J4i/Vq1ygXBHhR2kOJQi38WhpLGikG3vPFhRfw5DzlbIyuXCXAgDXYGaTVvtyp9/4rZtNT
GXinHB6g6CQ4X3Z9dnlhx2q70FdRfCRkzJQRDGT9EO8CMMGl7ObxKVjk/rvFKpPmDVtNSCVX2djz
mOndY8kncXP+Yf+TasxVX1xtsbwM1+Dpbrj2j+Y7dusL0+TSUBTE5cuE00nFGHivpI+wUJv9z47p
NdTIpYkMyoLKs9tZkuax2dVvV1UUgHZJt1fC0Ub1ifeLNCasMOnMckjwiPVo1RwxyYi/owaMPLZh
WQkKAR+C+QclFleoQpHP2P8nM8jMzRDesEArRiWeEI3DUvJq/dXmyEO0JjyLsDHSURVhaLmOIAmM
NtyPc8j6T54klQh3r+Mgz/Hhz9ll9ltEoU9ZRqmNo1q5Qlbh4tKcaGZ1CC2O5aTm1wXqzpqCBt35
N7MR4SEIm7jscH72N2bzzzTdd9RwMNNGed+y6NkiE4kvSO0UJxaBrw8YwMs1o6jqD/SE1UfnZeZB
TaDYp0Nww8F8EBXtA+TdlxxxC8mlgWtFhv4vqjniKJDOBBifPEU8/fNz4aHI+K005WjWsCrnHyGw
P8GyYOtC6GOlaRf2nI41JaJMvypZU5FwEs6rpyZw2Dx3ismgRu4+OguP+YPMHXr+WWhwH1mVJmUp
jAo5E+JGuv+GLPP5OHMfrH1lZ3f8Brkuiy/h1+Ufs/H3+c+BkzACvPbg56GM3E1QV6C52CTDtkfF
6Di5keYuZ7mjiCeEoTw/QIYpntr/RKsGwOerMwr24lLt9MPj0T6JiY3Ldyvv00LdsEaaI01gJMJt
/8PwoW1SoqL4DCVzI3HwX8pVk/vKIQnfhpoAv2MafAI7lMTH1v86M2CFJyntDs5ptB2vGp3M3zm0
WI6ZOPPEcLacrz7wPBL9mcE2e9nOy4/Fu2hZPOnm5bAbHD6QIJpxGxCobWHJ2XF9o1GKrow6TJ/U
dvzUkNT3FfnIgS+gLvhjH1b0Sqy34+1fUxOg8CIC7At4gR/ulXx5asQYk78GTGTq+//uFLBk6aXV
s1imkTGIqddHM/JgsqREHwV1tZFhidTIdUGFr2YiXgOrNTyFz32bZb9VsC0pon/QN8P+5wB/Uo3k
2u1TU5O5HtgXECUkxXCHIg1HuZ675/R1KNtJwtSbBH+DipKQ+4Kyg1DpRrOrswQMz9Lm05OLgL1G
B4g7qH2tzDFZuX6OpQ1ZLlSl1k88X/T5YnqbaPVoaXhAeM92yKXD1yAGbEoMcvz+SV8VJeirI4Ps
cirItQUzUjMTEZfIfOE3Rth7Yh2nCiNT3zkRzf75ZEoX+shVVLPZbVJtU7m9THKri+JFTcvrdi9E
AwN+wTsD3/v+T7sJVFEtTiE6HmnSIRF5idKoeeNmetGR5bzCeB9X8v/K+1GT8IN4FVpd87XwEum/
rztN6mpSsl3D/lnvxHduv/n8sHyPM1MgmeaHQpwfd+r0gj08R+ge2TMISF7llrdbvPTrVuOQDmZg
ZtoDjmyUvk+FttATAULaaM3TqGBjzXM0QEnO9oatoyuV1RGUQyqUu3p+wB1Y+58jniYPxy6m4OAh
/g0DGfU/ClMBIgXsMKVbdq23GmxtZXdYJpxkP4ukWMB47GRNuBhX+YHjCz6PaJJ0DztoMkjmlM3q
2zzMoZ0EB2FCiJuK/jpGnjH8wXdhM8SEiZWna0OTbD3yUz6ZF8/39XnlB8FjTULDhK21RGwl/OxX
qzIakIQA3iHGDfpHknAKjUnYn4KDzfibZPJQbUZeKpHFlyPpue5w+FrulkWcFBxW191615Nc24PQ
djvCRqYM2zoMdI2jx/yHSznWiyCqejZuUiPxXlliZYZ4156pRPkuMhY6usLbN4ItlCjdrqAA8Zcs
ebDT1nzAxOPEhiGbFagxEc2EXL7tuNNuVhHX/J8rU4g5FlIgENaNamyzCEcpBiRXY1bgEKqw5+8N
6p6YN9vnOYgjt0hJ4leFheB8JSriNOiYnjbtKV2bH44pamD1SykkUwD3NMSu4bhvYL1UOVblH3AV
GAnPbaSNxC/OPNpQcj7eYIidyFI/nckO4qWX+7eaBpXzBSA3rl9oaJF1MGyF2x3HVFR/iOlho39t
2JAEoYy7l01fLIKPckHDd+NPx0ulXB0+J4jJjMrNAlc8QGcQUscd0mjfTbST4OhZwAnPRdjd4DAF
bvtTwY+BGdT4GFwYEQg+w3FsaNAZrA9IV4+9gk5cLrPPR/6TssVFaajTGugD/3dWOSR50gxiLJ1Y
GQXrKp30mN3707RaaNdS0VOkiQIUFIk03kwb2W7K/MjfKcqfUPN7pf+0OCac3GUXPiYFGopQGtNh
AXxuMObUpZ98sIvXcAyiH2LmIOPa9ZDLb4vI2VT0dilcTqWXX/ywhgVPqPwoImqPs+HNPTpEOwaN
nmv5k7jEtYqnHbAqiCaNX8sQJ4j3rCLAAUyLiM5u8XSVsnYt3s6GVvd2557iswNDm4Eo8kQ3cMJM
3tKo6S38f1FxTlBVn7ebjbm52Ey2Eqph8HQ9kVn1bV9TXu9wXhmQ+wKdzYVBC0mRVMl3mmytjFpN
mx8vcIb+bakZsUd8lvdpLirnXfXhA9TlUhJCHKfBm8mDqtHmfl+sl7uQIwEv0CLA6YDb+kUZ/Y05
Lb7mYD9h7AGFqPKVXPGhA4SXucy7l4rwqiBVUWhSw/9YQIvayQdDz3r3hG2UPakr7wcpTPJmI7hq
1oaDKaEhFNe+52+x8ZNKw2GRXds2zeNSQJHOK6sopXCXOaTZKwePVdZ+aWhGoanJzYqdR/5Bik+u
ku5k+8Px08En7mM64VoKARbpH4j/IP/b65w5ICwgChmHHZr+Q0mtc6jO3Hf0aTTDE+S4VE3+hjO9
TCyffRLpM5iIv3cOydauU7yW9+IyC+EjDuCxNuS6A7e7tKF1OvvP6finMDv0WEyFE62RDI+gNEFz
xKd+YYnGrVr18tTKXj3uhbcmTARuAfwEOdh4VrhRsPnNCZ/YFKdNY+GBpMgp4f4NgOliMtlylSx+
Aa1CqWKNhAVJ3hBkS1RtCPkLSdFblvEctWCRf4odX0A/mQnPawG85iJVEQ2a5DkCO50XvvpZ+F86
OZUYxWBtdolGn56BvOitYXKAcT59CiCIyT+1aBC9WnBkcSu9E1wmpuG4r8npry1K00l1p+2eLcWQ
yLOBD1hbnYXrLfEwnFuMhWw3fGloyD/RZuqzfY/iRJJbWbqu+THu6OCjc1/OnZTa/+p+9u/P3ioR
SIuvR2vlOqp3S1jiukhDG0AEk1dfpnIVuZclaT776XhHvF3RJqguH8MbxVDh/wnrhTxYZiLb1c4D
CnmOIiOhwOpQL4RyoxVHFKd9vqLAZ7LTeaCTALROqbDnK43Gd+gyKa/MavbcsWKbkWNrOjjS/myp
FvU2KovH2UlWixeljqhnOMuJ4a71DuKn+sYpI9thC0XqZ24C3hSDrAshyn4qZUHky5A64kW9BDC8
8mVYfLIqzC7Mhtj+TcUzt2WbWRm35kI9PS3mA5Z4kaQzZb6nnSOoRGErIzJbnYZpkJcuz+C+D1Ow
DuVjx8QFQ/HqTsxxREQ0ssOE9Klkf4jdOsUVpgOY6jCpK8CFdRB68ENm0WtfHeII2c4X83qcfIR3
TUbcZ9A5CptMCwiNvKQnDB53BWXt2iMMciHt6/HakNrzbhZUzf3vkqt/3iE7lz4f5UMWEPccoKXK
g5e18dyZLEr7pOH3gbG6wkj0m7SKqrzcb+9x12BzOv7lb+H9QgK52rEtrQTKzvhTUJ3uJAr3CVpX
v57TVMfkDQTvurOYw7rNsPx4DjH27lJQZhilrQ8ftiaIt0hPS25Z4G4HZucsbzSqq1hkOOCiDgVq
Sa/3WCvAV2o/radP3R1aL4MK9PlXO9lpHWmtaz+kz9e7czDDyRROOaiy7ezQi8/x77l7Ood8F9DO
NAtfq9y8OkoB2QQhAGCzUg4lVhMqh2lsxfYI22gfyNV2epGuwL5RjET30N4h/VznIgtXkDYLLPlv
3wbPbIdjsLhJMX1oTyeyqq8ROb/FxnXefgvmg0vKfqm2iflJDKyj1kV9mhKNjSTEUNFiEoFcaJG0
MNnihYx1QjelS371UlX91MxTbmIC1nMfE5SJuW4nJHB6NclkTxsSh/N/D3CPoQltFKgurV8MDinW
rOgtCKiYoJXBP9ydsPknonvsktD2XXFszEeVAEy5busYOdpMnq2+4LtEHrtRtTN4HQ18Vh8M5oHd
8OSa/nO5aXml+xMaU371YweIxg29S0j8HfuQ0C85/JXayTqwD8e7zs7y4QYcvAHjVTYzOaZ9leNn
84ZLGHgsbQ0MAh7tYcgR+wYZoiv1gtvRtsbIuuZIAb71gLhkSWh6GbPP3/zUGl9lCUIsJwq+4hBs
T9/UY+nUispx+y++LFqOrW+AqOaq2xyikJcM7BuvK0ePkLgrDarY9ullYn5dMNaWRS2UcXxn7Mnq
cdVmKX07mLbyXyV6Z5wkd51RFCV9DLwJ/L/IAMmUf/erX5hDGF0q7IG3DeVxdRrzNRI0YtUjisLM
TQ4vzABq/T4Jc62PljQpXyk3SH7Dj4vjlYxTGUxJSYsg0Fmwwytc1Ecll5h40y8rS5jigbt+MXAc
q1Z3WtKqYjrymoiI6aB9Up69ZkYFS36ZGJSS79PRA5dpGXnCEzddn5lpcJpyNbswHAiaza8pE8R9
37KM/+VZp8eUmpGYhDOMukkQVelqXaNhOgNn3Lm+2GH0WHD+uPV5oRBCDS/FiXQUkc/iE47tz92d
WNY5Bhy7qzvxj6rEr+NATUIRje1Ygw+kMs9iYncgLLM8TfUIAdc33KnVVeKKjMcG9H36vOw/p2YS
dLAKBxrhb39niDkNQeHaqwHrVmPdjToBacvY75rBigl8tD/C8uvPIQg7Fedj22o7p1E6lBY0cY0F
F95KdQY2M27JBMNCf1aHyIS1OY8EJaJbm+JNQP6lynkj7l8s6EyE+zB1swePKl+4MJbo1awz5L2J
SpjIksPxAK3FcS3Ep48s3CzLy++8IMLiA1/7RprvR8UxSjlIQiYmuqxakCtjD+H8fUwJ7iI5LUde
uD+pecqfszS1WDGrv3WuB8Hi5TODzPi87AwJcVdxMWOwbqDdjvsWkfwvXl8KoK0Xcb1lGb2xG/7r
HDyGO2DorNmLZVDcG3ST4YjldrF24T7zypxETBG7N0UieQkOaBsRasf2GT8gF0ShmJV2+ZK5ZFBI
ySJ5Err7vJ247WVDt+etEdcOnUKE2a7kjia4JatljDPuEjTJAdzClZ8zKv5gW/nBkP7pSBZDx3kG
WasYDImtMl0Avb71C6Og/pMldobvUs2CFpof4fFBNk2sRPjbD7sc0H/9wmS9nw0RheCsixDnvrHF
D2nJHj8yFOcT3XgzAKfopa2O12lSbr2nLaFqTM5N3FdUD3XISciQ2egxKsmTfvERNMlGmsFq+L2J
r8yc+mQWQiHCIthB4rLzxOGWttfYhpeuvW9a9cbo99mv1fYXar3+uyCd/93Pwg017/BYGsVTYJgQ
Hda5OBJvItxclr93GjFkSW765/VF5mzEdGcVQhZK7vFD2brXxJwRQpXB+hTPo+fi1ZZq3Dm8iWFj
isWdtTyMwtbM55SYvcdAwjolaQRq3/J+9V3CuulMyXeT+H26Ud39LW/dZAFnGa80CVX5TBrAuH/9
GJWMznmFmTujl+nAZY4qKyQKNPGvdqtm83vzf4Cs4mX1wIT4ajd99RIPKs0bb1yKU7+7zNgFKI5Y
mfgtFki1n+LF02g0U/tWT6zrzH5qi5IvkwAJygW9k5bIAS36uFI4KeRMk+2+gtJRNtmkPbSRQ3lf
+/ELGn+4tyWWAryN83X5kfurUHS9gR7X28J77q8yBKptxxqtf8Z6oJBFTbCJhV2/RPf1r59O69U0
UYP41pD2pVNslfCyViXcWDzUiTGLuYCJL6wfEzOH550cSaQ89LeMUUyCtCAKPASKP3dMnwIesCUl
rqYyv1vFuYhxg1tJI1OWXissT5ZGkTM66PXs0tWg58jOjaQAqIVjhDiDqVJIDR8+ODrTSs+v9gyO
SdMoV7xpyVR1GR46LhFQ4u/edCkxl+B99f252C6eZ0x/c6qGyVcDK0wtTNpFjxxn/REBm6AxwFbF
11LExJnAbxBVlxbneDDrRxNRv+bHgfoHNsFotCAlRhszWk1yDK15U8MN6DGpniwuivt9m4+luLxL
9IihoreRlzcB01EcP8022miZi8BeD+QyBjyVw8vpmWwYi325wG2K0YR3CSOfDVnbyJfuMzfZxWEn
eUTUOXMdu5+pKS9cJ1jJudiVhLro62cYXA1sKhQWJVy/CeXHGCrE9S7uyC+fk0jMRn7vdnjbgIVc
JXMgp9tr9a7JmnOza1L5jRo6yNKVDAgdtuMyvlG0bjUi4wHTWUJq4kxSfUisjZr2vFuokGH8Y+qX
IrY5wxlfy8BMa3vLeQab5Qu6dJm78nRDQqehFSFPKJOXW9j3JP7GyZd0xd/TSywR0CViFIBpIjit
oBIpHHcbWzEtKIo6qF8bfjrfgUUD2ltdX7O26lJriVyOC3n6TdUE6OqxJNG9Ipr29CLRHlHZBc9F
AysAyqGiTHB4U0Ct6gHNgEdkdcWBsvkhQqRawTPBmQ6G6SFu6/byx5ohgGRUlOBCuEOyob9Fi75L
KSYfxKavlZ+vzSFAY2PMmSg/iBclMgWxlPcUxQORpR2ZTzb5xk7WBbiipCB3eGcCasZ+E0sqBbS5
iV+ASQzduxMw4dXZte2KTX3DOF2wN8IO1gadJKwACnolF58wtLs+JZYoQuuDFs4unYyT56k8KIzU
Cyo+ox+01YtQjWnfyYiM2vHWftfn/D6nZMbGK469zxHeAL+QuwJAnm5yVHDCOJMNdQfZ/c1y2BKq
x1G6XsVlqrEH37Gr3WWHXBdGHSCNAg/qShCgyAiYQEFzaSpciNRUIYiWvH0jU0hny1gyJRkUBNVI
DAMJhEPlPaTnzktxOBF24VbQdFrLv3NGPGTrke0HhmNQ4BQUFmzAl0NFSBeyBl/jokcR6k7p2Wms
U2Yd7BRfvllbjc7t7eyhjzUlSuq7Rd9DHqlAcQsxJ7+q6A0EP5mFmVN5+daMh8hq7vITLg5qeaaa
ZPJpWYR/jgljpB2u5RYLy9W7iwN9I2E95iVP3vlqatOVDMI8Bl4GTbBo3iX8H6063J100wLrwSB2
jwfMOetJZQTDckO6Sz7Hw5bc4+GRoHen9KQEP1IvGRjUABbuI4i8Mc1s406CfvV7TbOpjB7q72uZ
mxqfqhEMp0EqDiiuLGcXuJ6Pt2WPp/IQDHYkW3eflzWUmzstMw/4vin/B+ECAfAgKtxd+OwCfJT5
M5/VdhyembjYxO+j3JjvBnynOCWc4Nk+coL2jB4irygSQ6r1dE+RRcFVSB1qgNRAdnfU651eWPBv
yQOX5PK9Sgg5G5m6vkWpEKkT78Z6zLPejnPlV2uikrDZssefgXVlxFpZeBBvzzjZ1z+C8GB3O4AQ
DL5XKqZtP2XTN24KKYdd+nlp0Wsgx86XS8lgjqAbzuq92klYZjm7vGMpRGyGBUkHn1xfbE5giXjJ
wz88CO4ofskd7tnH8uOHoRqA/jLnfzi/XzA0lhBNUkifGiD+Vnc7AyG8e2nwkOBYyGex1l4SaApL
2c3c8Hcx89T/uItWZzwdQH7EzYVpjlkc4Vujtk5ermIX4j9Dm//vQAB3V6j/WjcKQjvKIVKvX3t/
y1HIkT3PYCbILQKGLplhldr+4Oe8eov3uHvxIhWGYzQhww5CxNsMVnEzxYLQazNc6zcqRqb5pX7c
fxMa7HQsP6Ha79ElRjCcuWCLL81X/O9HhDOTyqWqfhv2JpE4zX+4yNA6hwG6iyEeE5DsJW2R8MlP
TdAw2LtmxPPmvaMPSc26iEUqosxqFHF4hnhbjeQgI63VUJfCkhB9/4cjl/W8htddIUzBWZ57GXRK
J2OcPSacTphiBNv50KHKAIc16Y7mlBm9aI7v5mKJSWxxqbmCfdjSJ7nU+wCaOX7lx3RTxKtdrQq8
QXpJ0FzUEyHWCxmV551KV8Ud6eWAIAZ7wO05WNvqvPoffUXMpz7fnlB3BzZ84/yD3gnBI7YdouMK
A5eceJ7rzH8+PKKz3AS7Irhes5pN4E972cQdw9Be/2gpjlfYw/2i9xcCuq1vu9gU47WRreult7+K
2kJ50gHZgBoDTAhWqgDSH9jh0kN5Btk6rc5GEE0QhFYkWb9K+DwcKVUUjy0dgspJSAvdk9XIvmyn
nUX7kBUjPUkiUoxByQ0fQF8M+AFC3XT0AYFaTnSWBQgq3yGtycDetf8x8E7CE4igCMNlGjVDxLTY
n3cyKnPWVRBX52qvWe4I8SWoWZpjOLn82dyQj1bYBNL5LUyc/z09n2iLnH8tLvhFe8EntG8rXD1D
YXwBc8W/4hUk49Dq9S7RPSsnH7UQyNv3KEtVjdbX1zY+cuyLmnt1A11K/PdMB5cueEC0OgpluS1L
XAR0qmCXtraKGRMntrpx4r3G9TIMZxJzhn5ix1XURzcdvJ80P87xRTPa9ruv7XDE7NBrvVt6NwiE
dc++8lVjS+RLA4PG/aENecUxqnAmN3Wk03Bg9ln2wkaXMLw5vZnqMhtRwdL3fi6MPf0ih7nqGTxG
EkejQsSgpSsaYKorbhRwEND4ANno+DqSV6ktrAoCElOLnPwyGvwNADIouRXn0zhRWrlntpKo9q56
/2lPRZi6GooFFMQn95/WMx2T9W6kWHm05/fgLKg3Hzo5eNkO56b2BefSmT7WyLxzJrppA6xVaVhx
nVaGkrkdywWvZCls6CL5WrgNw9AvJj+mdac7EZd51AbZ2QYvnvGujvC3OBlWHsJ3K1E7Jp1MR7Ev
9kkQLlKu52SHhvv1Y6gAZsWUd4q7xuPW/Vo78f6ptyEXUVwMutZfOY7aelfq2VGzuaTtq/qCX+5C
vJX7a6b3/7a+fbz802cSWUupkuzP2PfvYJkOvQtNxor7sPNoit27GJ22BdMds8DWbtwyRL2zbdxi
WxVhUTmqKdx//nwraMIAmOptQ7iYg/d+EgJOi+xG/44O8L2OEzNIvgOiEqMV4AnwksVv/O2YVPQu
IjOvBMGwQtg4fKw8AfObHRelyiW5Zgmt0LP4r86QnSJ/hqyHsM9D26wKjohy6F2YLwWmDFh9Eivv
b5C8Aendoik1TDomtEwrLcrKkrY6JIGk98yY2qsl9WGTtxCfuayNKEramjO0Vn2ReUpEudTtZV30
b37XCJz2mixkmtcUtqndJPRItoKPeXnIj1v5szpyUqvhor9aLAE8KPJ26qvtS4LoiInjJ6ZQ0Yh2
jDJ3itCjnhiTGlpLtmgXO49HCz2BCsHZUWbPUg3ru/jJb+QY6tSGedwp7v+wfGKXAUz4A5tmHo6T
O3p7++fWfMU1YZifXsKpJfIBQ8+q63QeU9DoT8V3BYMZh1Ca9Lk4Igxtthbd6zzWNrmGz5vqzXYe
sPkC5g/hpOyDDTgllXOir1sQ/dbHOMhmvAPXx+Z4GXgvpPU7pUkO/qGQ81XbxluBtiJMqttj5h6E
MZPlrK4pdSi9tI2x/jUnszWW4GrnPYB6ENIVuhtelztMqX70oHxV1ryHub9ApkuaQ0OqBaS25coE
t2AY9AO8C8pqdn3OvDgTieQCJ/g6RFDmCJZOOgkPFTPL3hp6/Hoepi2odToa5qXnPcluiBpQXh14
9HIbOCumEiHs6q+EcEaeqPMrOJ11sRDowh9Bn1aXrcdFuK0cKA2L9DkgZ6RLufZUflCafuupvnIz
BfmoqmR3+IerN9VhN7Uh6iWWtfr2mbjSPPZZrdL88GaQq7F1jnGJOLM0lngSeIc4+8+YK8e7Dv2u
YnCwemnKqKtmDzpymVWsHYQ4V4uBe91UJNb6iHtyRR9t16qaO3mfoKuHzLspLg7MynY/cGqu1Pk3
VCRJYKU9sILsxlYUiSYciJKQT6jRnW77UuGJ0b9Qe+DJmYyiVV7XYNd+pIxpkloIOvpMSlahhaMU
Jn6Eyn7iGtZIRxtSq8e2IkSThbwvZpmoC4GhtvPr6EgPQ0SMcll44l88NxlXs29SWC4gmI7OGunz
DRIbLCnWMI1z8uh5F+djfXaj7+MxzWNTvkm59lQW2RrXIGdRX8ff02skP5jXp0YCD+sxbamDK6Hn
tW5NsRI/WH/ENYpYBCltpoRyNA/XPBEJJFrggxCLo6DBfFrlzXQ5HMBNp0snO2s553rK5zSjhcwX
BmyJXFmnwYMGSzs7dol0v8+aA/BYGyMjaH5tB00K7PSHQdVeyw9wgJ1+0+iBrnkVjbr/V9sbLat6
oJdvvwwBfts9l9t6WbR2iMCkCn5Du08I7imdUVy2g0GsCdhGzwmmWV4LFssZmmRcA1/623yvkrpq
FLWNpzvbS5VyLVEMesJZxCpMpa1DkNF86j6ilu1YT+BcpCvdABA64LlcLZaFwDmpKmLl6VWjEHam
Xx4H5V2EfzOFl/UUQKDe9p6aXbbfaObGz6oD68Bw6c+xhLQCF6xJJ+HKZbnh4wXfStErfbUcMYqL
mQHFZuvSXLzjVFyCoXRdu/qWRi9My7QmWLsvzVfFy1b78P122FK3LIAeDAmvzhXZPieNG8xKNEKD
GeWQcwgFAtXPwUJ+sf/wwisz/y1JmsOmTKSUGrx8Fnnyc3YEPxme71eKWWSgxhqM7LYJ6lezOIXf
qnOSPBzMl8LCBH8x7PGpFjtls8IJhQ6Wjk6YZT7+6jBb/jOUdbgc1MnK4lnSXr+pyvIpwoKi9yzJ
px0kiZLUOE+kft7BgANOUlMBGjTjVBskfCN1O/LdIbQp+p26HEBN2UjS/Ozt9wdgBGR2gTQs408n
ZMG2s5htrYPXEGUTewDDaCUkNZw7RJ8EoVPD+0U9KCyWJovoPgXHWEw1vcDSv+eJ8jH0uwUN9ZSB
LvpjAgbiezYxVJPdeAle853BrQaA2m+A6O1l6tFp2qYYOJuGlbtkHNDbqNZdbQqHYXDCN2WQtVm4
ES3ub2f7Ph/nW6+g3uiPhMjAHmyZXrCh3s8dm5S/1HE7cAIZIJftKgh81gaxngKwIKBTnROqJAt0
b2SBgubwc8bytmxascZ8aowqCp67uBnVHdfPpWxNiJ39W2QUjWRUkP94o61fXa/DrA7l/WpmQUCU
Fp197juv10CWK8occ7+t1aKmzP5k+vUlDFZQuz5coSEKlA2t5XmvbOORcmvR7zJ3hZOrV8NjtN0+
QyINDfin964EuGHs/d7OR5idKKnc1KCZvpRsWlwX6M5nFuO1OpokvjeIWrL3u6zdlmWUqcJMptre
H+85J4X5BlXWYZtwmahZqKwhsXJwat/aOaeP6dtwcnoeoD1iH+/HGgUBrWGPv3c632u0IY8dvuUP
u0gk2Rq/rba8koFzu0dcbp5oYWwYYjO7ctjnq3rGNEqC3i3Toe1FuBoDkDUt68fGsWPiXoEkXrCd
kgOW+80IUh1tXbsw1m8El4OkTwTqYDIshaAkGQofd1q9Eo+UcXsHHt7ypiCEzliDqSafrxBrNxb4
RmPdnzFG6TouTsnhuXDoe8YiTcWytH58XVN5I3hRhwCNteNtzf7WsxGayRHmgFBGdWyLf83L4WiD
YB8r1NN29CM17GXdw9O2K4p+nEXUW29+3IXJY3CAEFbjGqF6PTc//ycEuJy/nAmSST2dcou2hEU4
M9ZxNNO/4yBdPw3O/Z8HBoSwWN9xuDdCBecSxyYs9zT98El7yqSk7+H5+vj1tnaFYqP4yE/Hj0d1
b+VjbVeClqLg/0h2BYA4i752Taa2qzRYbT/uN2Vfir7hs4OFgR/VIjmeufDqk+/KkLS7ly4iw5r+
ZeETxd7vP2kL0SH3AgRrvFQqsEUZpCgKVG4vBFXuih3jhXF7a0VkYyWspP8OjhN6u4gaC3tw8lao
TaHizpul88DOlYfQuHLs1lsM2f8R5WFhQ0IrJBFhI+uh80qJ+cCBTgQxAbAhA4s9GfBWrmsW9sjV
IxVJrkZcHDg9ss2Lpai0M5ZdBcocFywufsuTrc2LAgEP6BgHq+1AYDU9D4QOEEmyem0sj/h4lK3F
oFOO9RwBR0wsYjnjEByDQfqOOOMORO35EaT0VCosJqEJhUEggwOZ7fVFiaBQsKijdzGFwCU20/CK
0q4xofr451vft7Iv4Dn8xoT9wEDgHAGawzdKqGXie+/XigKGfH0ekjbedkNV7lryfMOxoviIL66Y
TlvlxUDKsEW3uLpzAaMywKIO5BHGLYBXVxUW75T5E0gAZKkYuMctQup698zVH1Ag1XryWsj2RnI5
QvfsWnKz4clzDTL6J4hrrzZjTT7RmGXvY9CpUHrhjieBOknDlKTGBWJ4lPd4/j9VHhRp5VW+PxK9
FTosOlvaLYbAUN0PDLTtGzisiGe1axEcNd9UZFs3zPJEDtZjngNcKp1ZunfmGyuQiPcdmP4hISmK
jixKz9S8b1Fp6uiVqaHac2j9IRssxo9VrG+umcvkwuhzV/JhzFi/5a1/Obh3CzT/awgvlTZnJH4q
QCN6utwV2YcF6yYPWC/3rufrWucuvn0HfY4Gr5wqnBlPQT1bbjW0CzbcWz0pb5QN62LtUiXDmX8V
LLFMrYUJbvBX2no5Kru1/UKjbU5i7rfm6ifsZGzkc17VPcohFiNUoXWhzeB3WbJTS7JcKkMnS0Wh
XQnAs9+kmGDpOYYpiu3/GdAal8efMCvdskimnN0ZKEGt4HR19WpSreXD/hhpHr9/yC88Cn7jIsk6
05KUNi+MNgVyBw8x3cbKzPav7qm8je29QjwhmLm+X9lDnoVIF8rUxoGrXTkXCviBXtXQzN3fxtzR
mCKbpnqII9K9AI+DQV0W1/8IxsiaLXUwFxUfdmYx+cNXaAnDnkFDe7oi6X4ptOsVz8wha0/BiFnI
yUjojMtUtEFqlRMp5mN6sUG09rfxmRECqr0Ogg5JYaRtQWRIK1ooBxLbrcomnh+QuE66pkPHFr0u
QyFsS4LxNYAp4ckaGWlkRtaxHzukDUSvLy6D9lvJlxXuVOt6j3fi3ZTNqymZqyoP5omzncqqaIdo
W8NLm7c8LkpSN1A5IrQ9P9Sz8KFUmkol6/bSfpBK+SZFovQutTOYZA8BDX5d25qHQ50Q6K6cm5Z4
olc2OsrydRy2SAj9p+kHHLZRj3KxG9ODayAygBdLXsm0Ng69PIRpQQZGSwoe3neFQbiVTzD94U+/
kbEauj7quWznPtC/wEhHoN8/if42xE0nOzNCW8gYs0+08DU6kDaOPRkdx/+cu/3tAhWVl3oRY4oq
lLTyp0nvc7r84oNc6FcR2POq5Bo+WlBR3vcZTWtL+Ql5Zxc/pyMYjvWDe4kOQGuA/J9FOOxUahtF
FOe04fUtMkEH03l7Vozf+7SjG7QijqbMKkO2GW/ZyMS6NxzT5MmEQojVYy7aQY5y6PEmnDvdqJKw
z21MbTg49gqPL/doXDYH52DAg6SF5XPftu5a4zc9QuuWypcSiEcNG9jKlJIbzzQ1U4RXptwaXz5q
QNLMyixNaOsx+8R1FZ1H/9h71frjLVDjK6MCS0de6h0IKxT/2AkzjaU+nvz0S2uLviSHvoCgIeIp
hWdzCpsU4IMutNDqTv0Qq3SREKyaIkpEFxn2CBQMzh9b3h2pVNSg3LOesDpVoFuox2DczgIrn3hJ
DNG637AOgEgiD8uUR0qv+kWOjz2Oce/w+WesuLLBOJ96/JfJMvzKgDc7JsIy8T45TPtldY1FVVBJ
/qS5f3fpaUmcedavIUYLC5YJyE4cDaoiVe1ZKibQKqj3XHDr9pt9dCAiw2tf3INkK5wxVEz0Cmbk
lFsLmPJENW0igI/Iih4jY83wV/Q+TUANVK0wDueniishy46/1p+itKF1zDzvw+qihVCKPDmuS8dv
fVrDV6U4e37hzAZAHzhtFTQY21IMdbgcr+t6J1FOOVQSolnDafCB0T5crZOOqqn/7H095htJxD4V
bi9MaTriRJUPToQ9osOXV9j9KCxJmTJcvVEU25t9xUrKVkNAStEPNEwqzYAP+xhWUSsV7AajuUG9
612hj7H6Pqy6FOetChwmRNlKGy94h2VpYriekdXJ/IXfR/v/XK3uGGy3FYO7o8eNlzQ9edsAr3es
RqSK0LPWcfO8CEpXWmYm+SvHP6/PfdIG3eGQqUmVAFUrTaq76YhYeiqTFbfwBUN5ScgoQ2lSNwxz
6yhOPyWJBCu9wyfC0p9tWF9cF8PyNHqdOuEePTErO8814XI9MP57vnu+Ld79i7/vmxns7zLPQXe7
Fz3kQpACEiUSQFIDvD0cbF1OEUlWD5/OB01tdltwXZymtKahcBBGbNNIi0omRExT5YJ77k1DvlNR
WbMcHS7TDmBPAUQN9Qxox2zcOXMCiOQKcHq+zYEWuoQkM68DYxUqoLZSmwteR6x9wQXZdmZK/NRC
bkD9h2zzzWpW+3Dull0ic+wV/iNVkLS/o0OA/ncOHio/e+kuLtozGw7ZJwVt7v3SDy0LwzTiSVbi
VjCKNb8o4hLlJaxtcvMDiqBXTHVAyPNdBs869cqNfpdPQVF5rBNR3XE19UU90ZsVvTodXvIcuegb
fxA19DiltpBrFdlD/LFsFPsdfIuoIRJ7xK2B6RJSW39iSE35y7gtu4fSJxZmTdNhJy1rvsAysaBZ
LzWyKomI14vmk2XXMi8KQP4l+Kvzw8OZ3BCgEQ/sJ6nAsFMoFLDjmsc1jIUBwKHYY7EJQvT8+ziH
1JOJMZ6pVwQ7gZuWp/do+2zFWFhfuMdDivMKTn0Z/idT6aSSGe40dXWYOFquERvqSAXibmkBAEr3
fbwX6bLdRX7Qnm7eOaPkOOv4KBXjIZhbIyYesP8ONiU7Z7NdUInM6jMMB/m+UeWfDJVp2ojBD1z0
D6Hd/klB8N4IVXBBqCga3yzRZb1rj7vWJ/dzynPbe7a40SdHgEbFKAqxwFv3yRoxQKVCiFMgl4sa
R27vQaUcf2VtyRSL6VmzrpRvlgJVYDi88yL8DWemnuZyJYOIUV5mAqQsXtZtslP+x8PHMcLo/moG
HYZ8G9bVPpDOjMvzNqJqDfaQZFAmR+H8sEPobcdAGbnEqWFLQ6S7lmjypGY3vUA1J9WTc5Dj0vys
uhj3VlDTV4rbihveIYVsh7miyTXABc/k/Mz+Lw/FZmk7+qKT8RE/Mqn2WAu2NxtCKLe86oM05B4v
BAuQ2u52FDPpbwTHAVTt7yz4CEd4ChZ+fQwYXWXfOGpGPjBV0ooYmGHrNerzANsJQh+yjVH20cV9
lZUmzJo1G6ogflHy6ihdP3/Ie0f0Dn811ehZ/TIPWMsOum77zdyCbt6ta2eqWhJkM6eU/I47YyGP
erhWAWU7v71txByjdb6KIBe/gwybgFPghh5DqRNad1GLF0isr/WdRv1V+TNcTPHTtM2SOCNfYawY
MBsZpPO1jHnnVbrbtgFSC7i1QmGuVYt5XBBhYAIJVtnMGtyUeloukC1lnBfnkxmXzNivAZQ9ND9U
M7h2ALf+YmrCvCEbY1YtG0nMjwbXF4vF09f8myt2JhnW1GbJ5x0j21nLYlhIwJ1+bOyaadp+NVKO
2ny+dJAEMVt4DI8nQs/Dioo+ubGFgXiV+uDktcbaNPAqv+mg6MwGlyRbNBDf79h54G5Yfr9D8nWi
ddr1i7oC5YSXstYm03az91cIuTJdWaV9BUFkGWHLZApglRBAJX/il6W4+rLR5Dm/4sA1UcdIObzO
CrreQp13JRY2zU3jfjZtxXKFW6LyS7qLeZ3nE/m/w0KM6cIFAGNvTx3EHL0PDUiygcsDgV81cewd
Q2IMa2tTPM3nFXl8MMTqPwPW7BSc3zls7kHfsvo7IyAF7K+x/aPnlQ8P6I9vX4/GNfZLNH+7vNtZ
P531LqyLvEXVnWb2pbcznu//ulbzcmRQAb9cRkxRsEMO/Wk3Ry9b7FJA2eydw8XQbMfMh1ztc6nt
7Ajf4R1KcSynxLZJqlVSSCTr2gVQj8VqG9jPBGjSjOf7i2ua+dmp8AQDJ+9In3f3o0e2dSiuPdSG
mYs2+UX8inAu8gL49tF5K5bJcpYy4cc1r2EU7ijgAkjJ8oCOtwqCMPLtjcPK8doKAi6hy23NaW0O
VOTKAOwzqw3+sC+C6CXqhCa1RzmCZWz2aczuHiwna/Ufnf3O3PYLAmSOrFaOhLl2vFE7sFTsyAi2
nYsRBhcfmnRU7KhLWHc4S0nREz6yPqnwP6YRTGqJbKY6JRhDm65IEFuqP26CKyT/8lQym52kitgZ
Mh1jPsNjxBFpwrCKIYzKH22A91IdBMS+m0KDrfAVzWJLmJQH8h8T2W1XN50RkRohe687Mgta5vDg
wsXb0WGiosWp58ya8oQAIv1x/PCUK00r2vpMbb1L/afncQl4XwDnWFcxN8oyJJwgNsFadNLdlwKH
rT6kJwWGmOksvh5Kh6MdF51MhpmkznKiLqa3NH/iGZBgEHqOFEtW86xLSOztkT0pZpSQms4zwrsm
oB+4NWKNIwzCIq2mWnCPbnZ1uXeO5WaOxCVVMFyaOgfWe2W1YwXDeRoKp96InO24oNFvWV7TqjDd
gKoliOLvw6g6P314Hslkf9TeFHWZR/yrt2+W4fssxvRJYc6LJUtlXWV4IcsFKSLU6FXwSqtWRSM0
qlAiKkVHwozmA4cIjG+MhXJSRiIsA4MnIXXetPCnmNklMEKBlmyO7QEjUDgK/ZVouvB72wp7BUXk
uKWd8zjY8nEQsWuI8bt6d3ooYF+SJB6dUqBLGml4G2PhT2nmWc2Oy6XweWPa6A+IDUMZZqDtCLuY
2HWgpbfUnrklLwU9/u5PoUaMhOoHrjo0S3QHsxTG16yCBPE/dsoKMj88pV5VyEBf9dU7VtbYtWef
K4fpuQQTwscCgjjCY9ZGv3N/IE4WFyCCalg5gdPfSM0k5xhIMFGmeD7BbNtVBVT1MuzZ+nREGE/3
ou3UA+L+LeHh6x2JpPh/A8EQPnJ7xseL5UJrx0JCLqAX6RnToep6av3//2BVKy9/aVyXsgQJzOaA
w8+YK2XxKyMkieSLaUJo6CfEfqF/do3ra1e6QMWmTiwq8fnQ/Xb50Se3hn7BbdNX8M5PHBX7ak5O
exkYqvm7cf3GOmCc6BkTiAaK93ZYxBGNp63MxdVPUWsX900VOKQxZ6EEvo5Ldw1jwdvL+8Rp3ehI
koaLqKlJUd2h1ECsnVyZQvD4+CBoWHZV7quQjNvrMiT8HfPvXDD5eT9TCOXMKqXO+uJY1uUZsHuA
ay4B0QY/k15fwsPdRGI9fENfba929p311qu0pd4JuF4rhgprGx11qLHut9Qr7N8N2adXAzJ/Qrv0
iYLYguXQGB2QxM6jX2k7CfOFjN8e8RqbWPAVm16Mzwu9DCubnVxb3Y0Qee0IZpObIgrmBokg0PxC
ymLw6IBkvHYUiqwPHNp80yKD9cHAnv3jAwLxVgd00I+O9gl2xSPaABIF7MDV7OId/cCdv2iDvL+f
1koWggcO2XUv0S+5L194O6QZVl9mvT4KRj8Ez0qMjJ0UY6kiWvF4P5vx+lhZR0eErSR8aHKr8g/w
TuTrysCU5UHd+SBWWFFDPlDS/pJkzTvW29l/om2pGgU3sYiNBX7auTUJs2KBEkdGD5GyffhCsJb2
kQhuE3As+UfYD/r41HDC4DUpZDL99mFSifbBL5Auj4SoOcod1X5VKq3PdDPHKvgpHJGpN1tjLqzU
Tu7xxTpraV9ATiIARYjx71eI18MJKRLAR8sHEJrq2R53rmYBQFSbpgtS7lDfI/XvHdPKd/uS50AF
MWOnwsGax9x/Kz0EgCWJTTsFiijvoOkQaJU6nL8C/oNA9CvdqGKMBmtvn29AyAGAL3luiQDf46HF
rC4jv4KECQmoHeRS5aTqv4qtWTdtR/3Y8FE2tMl3YIxE17CvLe6gd8GOEo4vWdgLbG7vFX5bXd4x
FsZwcvBFoJcCcI0fJL+QHpY+7Zcsa0Ezrf1FhNw82+1bK4wgz51zVgze4HnH5OY3oji+VZi7UoTn
dVG9EZQfUy9HD82x1Y8UwsbtIAFu5PzYjJekCEcQZX9r89fmNU8f79Ko+6/vhrd9gl7TYRTNa/fV
tcHe8075e4iC2l/hVhpdyKd0nDD6n4m8iFqLNhDGs7/Fr9+2ocH8HF+/vbgq1tz55UbRQwUj9Np1
F43A8ncOnNVhtX/tak5vWK7qXMsljoJ730bC1DxPDOT9PyAix3LRzDmlGTSFMUBGdJTeWsXZ/jLU
MUIGwYy7e2Juxegc6Gy+xCqxmDB330/2+AOd0WZz2ZZZfVTUlkcprLZgo9zcgLFdsfY4bOKmTsCk
XxHj+C1oIpcsqLyZs8Pn2rvUMx4iTiDxzsY37WD+u+7G5wXb/+ldwnvPRrisMI9Wm/t/AxrNtg3G
+Bn89Zw2blT1aylfjYxAtStjSxgDG5A28u4vHMHWle1kyY+zpOV5ULAKuIIXbmgjrVFa1TTYwfQc
1w8tq7L1f6RhRT57DLdncZthrQ/pEuMBoxJfUAfxAW4IbC/1rdS5xBNruWzkU8mcFjwd1iJ+YMFJ
44rxnGL6QAJJgcgA0Hzhb+w3tNvocMhCSIScyfPi6mSciqzRgtgaUpTN7oNh1RP2ZQLZbczAvo3y
IGv2OidIfkXbInkkwFcWRJQMLquN2ERfWMRBzY3WL13frP9v56ERio+2vaMs5EcIc/99zRJjn92A
vAlUvVuTNJCONT564XpYJLT4JsFywKpAGlpZwEsESplvSY4KLReH/GMQxB3vWUj+Qxzda71FoXXC
RAKCq/Il9AgXybZQVtnOyG7i/unmcsaT7BLTYen7UyKL+59MlWhFcoGAxm/NfgjIfmADvm+2tLEj
SnVhdiwKgxwKhctZy3HeK9iWjkdnC/TjYjR8V+/PRjsa8//qCE9Fg5JK/ZW7GVOPY/RjrshWbKqE
ZFnmgosWwEAmeHhexpkASNUqNZZqZekFK65GfEBIx7QVmCGgmxtga36rTeOKTWeWalur/MOMNaRF
6/vamzOacy++tqWsjyiwpMRcWmSu63HD6aKOZV+RPUM4otywc3G3W0jln34NBGILwmwlEhHlxGSh
+uXZDWSsGbspCP22xQOT37PTUyKylRIu+z36v16wcVmm34dzMs2zhkf4haMSPMnWG5zUy+O86Lxw
d5SeN7JydXH6m3Qk3Jo9MEVmGhw12QOROMMBkoSdfx+YG3rc49KQvUzk8UA2w9jCkr1+6Daf5WH8
MRTNdrtBT1ZYiXAyhPnojp+12S0okP261T5faIwdFI8aP3vnnfXeVA72iPFx07OlX9WipcxPLZCQ
QT2Fvznx9OGoAaKYcHO4y0u0JFS41k63L9Rik44KrdLaDZ1jndx2fVLteopiC9KhTLECIxYdF5eH
tDINry+CrCNwOMlkdPtMpT7ZMZUxyISNugICL1AbgWgDlY/LE31GbtwL2NdxQaqAGpRIp77bPjkw
TOr/YStHoHyvp6/qFKYXRbVfw8qake0BhUPM6GYgo6pFTnt6jL9uT9m3jJxeqLvd0NWGKytPNKEz
JbWPqUXK3zjZG+DK7gyv/wbtJnEJfUsWOq+nF7veuUKb9+bNWyhMCN4mRltHlw0AwDSSJTKO6Cks
bioWUvar+sXL3WBUjugc3+xz4pQVfISD5YxHhQOWHOX+0U+Tp+1LBtjmew9gaA8lhx2bojtukXSs
Vh2NO915KH3TaR4zyeRQL6FH9SklngJhwiAAn64PYaMZ2qyhylbQ6dWNGT12+ab7czmYwffQiAkJ
K8fAcsOR1MOUj3qTr2fjC3eiKEEBbzp/mkU6sUvdGPBKTLHR9Rfep77lI4PIEAPcMWa34rkut4AE
YixvxX7nwazPnAGXb9SK2LnBlgovFDTI3DEpEJb25GtEgDocE42KaJ7IGkntg+rVILlQ5GJZjS1y
ie8kbPuh6u9x6IZkGLyRZhrtsRJ3EFr8He5meTuvcKozc4ZjZZlQRH8Bl2r6Q/gMa3wks1yfL4nC
Yu0He9iIopIbdILuRnMVypCk3r5cPNlq6SabaMs48RF39Mx7BHipLcjVasBMO8z8dU8JeAUKEBUV
f899bX1TcaMC3CNFOObjNq4Ky1KZgEidN1lyh0y2NnIKEg7LQoznta5ub5li4pnqn3i9VFYhfpVF
PcYXkuOkJW1gULAiLkPXq+/q/F/tYRWL9ODfeKKdsM8nW25v99+h+AiHk1r5nQMKHnQ8Dv5hr1nz
AD4tZat5UFl7IubHsFdc2d9lyRIKp+sj8t2RNLMT3GlG6a87CbkFv68nNjN8H0opT8GY7lcR1mfQ
mfLF+VHxyvNu8kXZaSBCJyEuPvq/fy7Moc+pbUR+dBPHIWHM/r04MHJJ7tWe70fqvNxr4b3zD9I1
a6VvnnbHGT609eO2VkEdhqhBM+SNm+D6vqzntNWZluptpHvBps6m+Im4D3uxnBSF3DX6aKPSM85i
LeUtfU5qS4fFKsBsVzeengyIRDJ3cNnV1N6GT24BibPq13zurXhmOvv7olPx3iBvhl4pcl+Go7DZ
yGvfpLM1yUaXWf3W+iJjyBRBvUiwAj+6aqejT8hw5sauCF7N8a2G2iGpMf6wDW52S9HBhazcEIto
NB39kVYcMYQujbv7NKZuSbd4Aua3QsbWx5drWXQHLH8MFN4mSHZnSJKv/KBchz4v5MxAWORuRCvP
gYiA2Wjfvp+nP1+Ae3Zu3E6OWP7fCQ9ynyzy+szS2bhOH/AdxBd62aJG7hqbyN0TITfMSezax/1o
cLsqXIIn+ch4ErfMUDSzHGpqtcU2TRFUerhIzft81BNa14g7v9JZWYCFqFeRQfuPjoPVgBcxqZhm
CYt7DFv0cwKJS3WxwhZb/QyVJqIh6r1/oLyHgABzInoBUGsrkap28x5mMaDiMAGSZesqnddZpR34
XdYwjiMcor4DIQ1G0vQ95e5Cs6/VTK6SSmGMT6y4EubWThAau/DX+ADCUzIrVT/kNw23RomXNLG3
2Ruw92zhtvjww+4yPh17D6ojK7GZjHqG7Oyf7uFOl+3AgYR+1kQC3ogJ+ScsXGygb72UqvP5j8LP
JAv2s0q5grfAnSMnWoY2QDdBWsC4ehMtcBmavOXuLoapA8KsuH7tQWZFoxbz6cQ61G3WKEjL6Ekl
9n4adDL4utML30xVraf/mP+OKj8JGzkW0dzI3/NZb7FGK0Hev3GiE2+YRNkPs9EcElE3Qw7wzesh
wFIvYWTp6WrX06oTEOgQP+Ocxg2a7LuBCBfwaVn/O+5JKqDwsYYQ9Ne+4QrRt1tvtHTUh4I8vGDx
5sUwkRu0jS0obeDGRBhkKgG3E4TbepJisux4q76EVjyIt/PN98N+A8fo7LSz0TFDP7sv/TRH4CpG
ur99SaohiMPXXZZnKCZI2OXHxu4ul8rmqPBUaAqFp/SftO24nMZTaq3/DIZw6r05VLk+Ux2fQy1Z
F6D3wIxuMf/XE9SHRH33GVH0BYH1Wtp5ZpdUKXaU0gH2JI1MSznJjf0X2eMiDAidfXevTrScFcn/
W72KnCUPUsXYQ8AemjLqQFNezuuuXdIeC9BtnYxRSIo9BFyaPtcSkaHMPp1cwZkQJOW/LywW+8vT
2dR8WbNbcRxkstIwEjZ9f5cHRQi+uywU9zZBHWLT9xb66eFS46H7mKW1xxZbXLE+yw2N0ijdpPpa
xiBm+iRolUNuNa/i7iHuzbOjyOezvVnh/lg/phyghmR0absz3H01OFw1s25jk2nzertYp2EcL78W
N+Cgb/fYjYfoi6nlkaQ4yczpcJ8Yuz5T5MSY0PExphTl1+vhlygW+OrUOTB2wvgyg3a/+sc1lSWG
UpGAC+fa2CAf0TgrRvX1ACbKdUoxzakeTz/gsxWvjEufoW+O6vDpYjFCDU2qOnbFgkbrIITChFEw
ODFBxrtPjy4iGCO5Ket7a4n6gCKA/2xUdqPadt6u4yL4vsnyROigNCu9NB9LwEkYa2gW5OHD4FEh
tEIDDsXoXBxTRAC597dkcM3JWMAo9+L+q29Az7QN5omX/mBiWljYhXlVVF/W9RqXqwXafliLjN8g
Z/lH/R9pMkFt27Fz7cRGpdbow/VHO+5JdBsnzE6PBhnJDK1SDPijq7QyxQKxI6pd4R7s0QdZ43dL
KJlV/WACptXTIZXMn56I8kIeKveHDd6MBBp3JJaM0dWQPuPg80qnP3L3tp3JUhBykOVdorfZjB1k
GXJ+ZeJgMYlhjOwKvJcGqtPH8kAgj0BQ3RLst3ujOLPNog5YrJ63a9u0qSGDL2a7clJ64wjvkztX
hITUZWdClAbK0P5eYN0i4vNSWeC7jz38GwRTgLVGTbXGT0+LPOmGKKyYJCVI+zhJ6QCbAg3gy2Ct
Hl4z8b+MiLX1HfHJJHDPPi9bzuQZYt4Um7r41QMovbELWWCiQylNoJiOt6+ZOT9V0AqtLvdfOA0v
kTuDWIn7AfhYRkZQnKrEX/TdBQSLIS1gMAapGf3k8Erz4UeZPRiooHZj/gpRO/5jw1wAirr/oaHv
JBNGX7kW19b/c9VS1M4QQSE+w2fSIh+Qc5hg2j60jgJWgqbpeastEXbFLk1mnhBVQMAOIUHxdQ4n
3VBUCXmugbBkgPhcBLcuUlon0X5rZsDg3Q4uktN2OnjjcJ4wVAf8IwS+8h5UVnsphtJ8RYee+4Ii
scfaGiGY78+2iQMVhdeAMaitiGvb2fB6qJCRCRuQ1lb3y+cVwJ6tSiTfTbQxq4e0uB5ONNmQwx3o
b9CAolvEySopmZjIy7taTL3g7WzSa5wuLTfZk21zD9z14KPiK7hGI8o+bklSFVIDivw2sHHaPUJs
7jpynw8weqo9w8C71DP2IpV7v4Mij6dXNV4hrcgmQNv4laHH3zsD8AUNMOfJl30wjU+aAGVjXOIG
MUUIsiG6eZz2CJnOAANUnNNEJU+RvNpyI5dU5qtb9no3ebdbtqB8Od7lTzrlxmwnYND+SZp8zHHo
W6bhBi7IP116IW8hAuxyBECxsemnTuto08Bwkoz4kvoH4YhYXt08upYsKATQrMZL0Mm56VjNy8s4
Krund+0pYIBY3Jy/Mb8K5Xz9OWMDX3UDut0WSkcl+kX/pbPEroLeujMjxT0tQPTrI5qHty78aONC
J5+86qa9Jn4bRbgpN2g/d2vWCciDAnpPb3/XaTX+PjlVWPr9Ox14mIQxVSrF9xL6eiQ1cYkr5NFM
to+ABVu/MaHcd9Nwxv9o1kiq4viplnTE3oh1i+6QaNHI5vTR/+SrJ2sK9mEauzRQ7rETwsN1MkDe
F+CPYpZRY6USMpoCjVLjGjMYzlNb2NQjFih9+uhckepJE3YsVxB672DHvNxOwLJ1HhtZsD8Ar1qR
joun722HK5KD7Wi7v33kPu9/hi8U8mKyoXjcgbOX58OjMxZyGk+sOU6Hp1l9LxC4h0IIEq6WTG+a
f06aQ+HsSrI/BYayPv/eeuqz6pbHVGGYXhawCGjhK5S1KajfmeqThSkZppDFxN/zCu/iORMDRXJh
OohwPP/sbjeXyUroVdIHJf+xTcQwFtJ7kOi0srx98gbaRugSMC5nSy/0Zj6lVggn3943QSBb/SYd
Ne5Q8yUQIww6sL4TPLGxtrqFYrge0j113i2LS9FLFYHNeA+sod93lMMkbeSaU9PlqRWOluR8GkcK
ficB01gowbOKy0MR8QQVjTQWLjhBgfbMc76yqgwS6qB3AJVnJzcwGUuP18fd1yUjYSrux8RMXMy9
WSZgqDlTOA3bcSgOyZ+374U12poJHYLe3/jkyzNxSc1829z7yRwSQigD+6VILQp7vESx6uDHBQ8V
wX/JUpTkrkCSi4hbfdsnAjG8ldthysXsxXW5DikoIgX5TOBZk7o1txjhptImRdM5Qsy4R2wIyF7Q
k7QbLwQjPVms+Y1d7wf7v5AsikG5EBNr+wpNuNu2OotxY+DL0EQblj5SE8CnNJj0oMdP6QeyFa+H
/eyBfX1pBJpHO8lqmDvq9acKnqj/hjJZEvwaJH7uE/tMLkR0iAvpnXi0hqHDJQkH7Qdpszw6y2Xf
wIP/TV8W8kM8xQjkKrRcOYcLRmBmJLVBBrw1X45NBtGuOwVcX+/2ahORhrEGHFrr++Pube+IRkkV
/A6pIZJ8jtG3ugBKKDcEhRi/SCUFo45xjQW4xaYdupj2QD52JjVL2QL3CSI9hqGV8I8T6Mqia+Z0
Nj/XmbWXJzdPet9ZTTe+vU6E8dt2/DPj0o6ZtGPU/E1o1ozp0mMKZWbvxWv/BxoZ5SMlYGAbh9kK
jA7Lwbs/rCUR3Wh6Yv6BW0vH9Lpq2PupUtI1zNQiVoB/3ULV8Gn/yepbh5kbqZfdYO/5EHvaJray
fR76u8y0OFvcBjQKQF2iV8A4bIWulHPRN+/0VNx/BN0F4ufBQ6C3h7JZ8OlOFI8P3b8fQs2+cUNF
EOmnOsVjcLBsaXmNwc6ADB1NWx/CYRRtjZqzsYzNvzKiUNWeJ/HpbbUOOSa60c8iLqyJ+1PsKckN
Ru0SX7/uXP/CHkYqzEBhLx06CMnXsmSSE6cgFcJpkQRz9STKNDLSrUxwiGKEXmklkbJLOTrlOXJa
uJZ/YBLAOaOqoizOGNcLaZFuXFAYzI2aSbouDZGNZfTsPYXSyNjcLf1DYn8CucTDPfwmwuvOysSS
EQRuFGPxvjoa2eD+YiLfa4VugwCjqQW8TnEN82orGH8gdowXjHMaTeMOqoS36Qtr7ZmvYEhEEs6s
tDS5Ou6sbNTQBOjDnJrxy6C+vyEO/6zfEVnt8Xusat+OuEFC93lOY6K5ycjdBQlBARSQ0IRU/zS2
QRxmfNKmvwlOzOjGUfCL41BAmgqwSnJsQ04Sl4AXdMh9jSoTN3iKDUYs8bvw6iZWK1QEek0yLRtJ
vyoPn0PWu0iFhIL6DFvgpLn569Q+COdkJnw8/w/ZjB4z4hjLjkQnQvZPOoe8Mb8ocEVAw4XfU6dD
l4HBoup/pAaFk28wV2CHV0ImmvqIQBClc7at+XBfvozcQOyDMoWbsn/DY0fSCUfb+wwQ4hQd0whl
acjtUPfjyr7N+pU8FOFURwECAcUD3YBH1PtWsQ9nWq4Mn9JTq65SL09rwtWAM9CYC8mV6who1Rhm
oAmSNTT6Psa+WyHpciNAF3pY6B4DGHKs+13nEvVgsPoqCgXg/Xctes5lqa5LtBv4lWU6T+2utlX8
3wEB5ywQGYoSiCIPjXjIGQz1dl86fJ1WpCK1t0kmdRpqP/3wdA4CYMe/7iIYd+UWGUlNIwQe4GvT
UTs5rpmp+NKotB3LjaIm61yKuxHBtgyvkoI5jF7mBvccz0wi1kwkJKxEpc3SrSA20jebo6Y6oI5i
wzA9y0h3pfmPBmSDyaClDC3BiDOW0s98BaVKCHO25hDw8fsoavG21mvJ5D/nfGEttGmmk2wVYrqu
EcB4HTzp9kCbuXNKpnOYJhoIXmJFWQjzpSgn7QbzFVttCzxkhqp1dEnhfOavToJwOLGX60fQ9ZpB
0siopqmVoTGq4znuYQN3vG/sFGh1R8d/ZvFkYIO+KwtiAr69/+j1MgGMCK4vC3qCeZqE9DNnEL0p
HRbXD2G5XxAmW0am8KbzyeUb2tvLyd5IZX/qtI1F9YBwogyJwT8Mr1Ms4/ZeThC/Tty8TS0XZmel
yVKmnA+HhciT4AJdWZiTYWihJT9bYTf55C1j6W/NEIeWA/7oaDTbcY3KoN0RDVICrgWfhKvxALbS
VokxWYKHTDo44TdTVJLP5kCb1lp46hnLEaKGzp0UFDfXHpjz+IH4B1VYRn/n+eyuBg1/+/WC318r
8+wz4O1SDwpIv/L25CErzSmbXBNmSQDWw6UysbvYZzMGL7WRA4ongzll1ehF5Aozh0Oy+wFDtsc4
psZhHqvoCVg33hw9CwXi/qZJZ+sME/y0qbf5+YdAKhhQeOPSoYhAcV7Rz7ul+N3pp7/jt2xK76C/
kVwj1qYpN/YxToh45GKOYqztDeJUhurHeD5YxAR6NuuolFNBiy7+wTUMww1Z6nounE61bUtbAjQ6
KHGArq70dhLTXZdOWcBHl8SDyD4QIM/IEUBTnbnYc7q8Ae2c3BqP1npKPY3Aiq+Ho6t5C3eUgv41
toen6JFW7lNoyKbd2rZoRDONyr8hEt/evWo3/92fkXqcL64c5X9/ksW9cWWwCPycfUO9AUIgcQ+r
jVhbGkSVupQ1FqJNONLPNp1BER3EI4PZF8ondWnuFClnUc64yja+dxj56Gac+RC+zTJx+4j22xXg
Ec2aUz5rbJqLn7yYwL6QoCZWUOdivXSAbyq3DdmTP1DzW4k3j11WYHr0YPvuGvaTEycOqGfthRGb
HOR4BuscAeEtffQ3H4oCJnHGjQkzC2NVgK6foffU/L9WFbZPRYk3sta1y8myChM+2Os1wvKD2cb6
suZQhn4samq/0M8qlJR4s8SO3NxD2szwwSPu/odSguI//HBM3NQ0aumT05k+Xsb1RSK6EmCICouJ
F4sY0DkCUqnvXTmmpp1o3lvGVtPa+9kC1F2JOT/oiuHZpQJUYLJeR60n0rGpLOJnKfeSMFZ+eOPw
mqkrLhKhmfWywQ7mwvMrO4mtEtt+beLpEYKDYBzCwKzsC7Ajnfh59veOS/FbIPR/uTY5GnlFtJOM
8ehm9zcxreKiIfzGaXm5ytQY8Du2e2Bu63uOPml6QUYmZiqJ/NZqUpKQzKANLA5f6j7jKiJyE/hK
R5k5MReeWIG2CSVxb56GPOpcWclur3d7QaSHHzr0VnoJ7HRWHDYHHm9gqnllkc54nmk0lcZPqTkW
pbNbPStlFOZyggFSDSVwNPMeHL8xGqYU0d60E/nHatU8+RLvLergcjh/pZiVD+uC+DNC4d3f2Acf
aDHs2CYm7NNOUw2qI1MgVytpGA5QDw+oZcQjiq9UNJfO+m2ZlWn97cUcUvZ2q8qOQ/8CNyKhsvNu
tlM3PBvRP6rVGBb/XJ4jjRyVXpOueRU2paQW2/RlShlrzMFJFxMOBdjPKmiaHCLsxvd3yN0z9ZrT
F8xC+Em4RqgflhBrSIixUcBRQSWNAKk+7sYZY0DrHgatoFjzqipseJ+EvhOpCd/N8W52XS/giPg4
fMaYsfhHlO4mswJkI5O6js4wTug3263ARHbILgijOZYNaw4zH7CuoO3YCGlpHY7pfYkJrD91rqhb
CntCXVbJE457YoVznbCPlafsBhQ0+dUHAal48wiyoQxS572sVk+k9nU+Q3d0phXPN1W5SEX0+/P1
IA61F5puQQ9fA34v32rDBORZPo2Bhh/dc16wAG/HKyPoEQ19zOeDWu6jxou34zxT6xBARy/jtUWT
xt5NtlZoQxpsKA43hEz6ieV53brZdiy0NaWEDlTNocQMYmnnYmGcJlNtEBob+SShnfQWcmUAjKZY
4XED1uR7ybGTXiQgguaOEmQ+CTQX+9T7Yv0j8HkqwbO2LXUMqWbGh01S9VMw8ii/iI1Lq59NY07h
8R2CGGW5aleUXTqQ4mqOWdhYzG81rArtUCzpBrEOZDpLbu1Rpk7+/pC8W1k2l0Ssh4ZXKmZRx8q9
cKOmd2aXgR12mLBgljy+r2mY6NoAVGRO8gGI4N1teECnAUoLD7CSVHfbgXTs5doT7TWGs4kVDlj7
t9tqC8tSPto1J3St2/DfAo6Y9X/6ocmI9ZM3RSC1Rr0P6VJNY/bskfgFbh0FxFaynmwgyVqCf3oq
BIc7Hpmx2Ex14t6ZlGrOLTD+EwN7pmlt9MwjubBoi2PzEGIYRs+8jnocqLOD4KlAVopxGH9ElMOY
gdNEbTG078i3AAGzNRhmjnY/RIklOwBe7OUyMRTRyuvZqCxSJudQFwM/DAkDGzpIf5w5nexOW8Zr
2Ke8/fqux29JwgTWqD/8S6K1g50z8fQ8ZUBCCSa2t8DzSlw/Tq0SrKcZyzM50fdH2mldtMdypyJ0
QMX8TC7IewssV3P0HRfafwMgSatj9VpuFPwvYUh6LugniV/lVXsJQ+zTIgyMT9pNNkXr52V3aeo8
1gcOvmPwKMds/KzcnU5/Q1TRxTh1HvmL2eBSTMS+a3IkYmrkb/pPqF8if4uOccRdkw8wiNgOsh+T
FxvDlnujuP7larlZZgdsZHld6x6pu7oJHtDLkbNF2A3yWjV0hx3i4g+FJd6qdcqvPGKfbDK0pH//
D1KLvH9lEczaEm8PS5nXndoqe0lzhoqzi+JTiAibpT/6wRyyyix42kushD8HLzN7IKy+LV4itrwp
QIfbNRRxs2VM5XjIgbN+Y/m/UkMHvzQ2ELqJTxFxsGeB1/5G/ywW7Eivqr7tnye8ELaKdj84jKTw
205GlvWNIRANZN42TUCfVsOiK3s6PG++Hcetci+xaOaHWS68nZOGuT4JJGdsupvoLxy7XpBNRYux
ZV0gGPR0I8zLDwMW9hO6lot8kpOzLdWVidWdFijtCF7IZeRZZ9r4bvC3/O3Tka/OK7QOQOWPGnq0
ZeQyZtv1blPnxJvOA3ldDndRcobkB68ajhlbT3Td1HOV1diB/W6LnsmySYInC5B0r3H3qWKWUCJj
BzsQI0+si0HLnYv0jX/Tf16jyhx2SDUx4GKG6jtFeRxvwlaFKdByqgfe/j62Br1K//zBjsPmAqQM
3jHfVQnVWdpUqjyzHXoY8FJz06kIQoLlxT606a8Fv6O4Sn2iOuBF+vtgGPTDOXaP8s6saKax06A7
Vi8J2euGOqClzIFikaKxXwdhniHkFG+AaZH6AdQdKYBpyr8rtYMSb3O8unx6Y/sd/t0BTqP5hHiC
yt6OWNoZ/uAbDZoNo0Jj1li67O3hYOEFeKtqTXpfTPPUw3cy3l8xoD/MqKObppM7yWdwa4TBt96h
xEDDaur2TyP7Kci7J86eM/HxHLG6N+T30LM8YgpfvCzxUWd5WJbGg7Qsf+mLJApH0L2yoLHAgt/U
8pIh7CGvYIWbuHVh8Ab1ZaDhVeGCHw+EUCqVbzRs/wQ2t9BTEiaNVTXzZ/pU1Ybp1Q4OIG1883SX
FV+mlACf/wYzug1K27zpWNyOorhk2x3d9C6RuXo5HMdGBrjxin5P0derdhmaSAHEg6xm8w2a9EjP
wlIOBITlv3tMcqO2v3wNr+xKDtVqxGp84ewXqJ9KL2TsT/N9BKPP9XxB2ZYPQwdgbgm28rcE4diR
VZAD6YkkGlfPNgYVcSGkSkhIhq9KbdR9laa47TAIqJhUOboC8jqKCESNV2yW9LK/Obu0RNl6M5EE
HoGxGZqlmIP2d6VrKoR7FfVuQDLarU67sLZ7U/9tMP0DaA+2wdcl6qINgZfl0pzNl7p7sJx80pMo
TGSsCNWh2TqYILV5DAeEYZArB8L+/mcuj/YakBwyJZY0SzjaLRaaInIO4Dm4WyMTPyvU8iULWc5D
iRGBcqQJ9TxX0bVvC+5TxwarMUHj3E/N3xvCXiHahfLK4NpWZzp6JRqQAKUBsS9bTHtz+X0U2TRl
5L62BLUohxFKuGgAJu4r8OiK1yurNwuFpdcaxPNxbY1FxSEg6uTtxjEXTKL7Z3Fn93gVlfNOGl+o
KwFR0Iu9oxb77VeCPO1f79sJ5kD912EUE4ViJwDzBW0AC993IkfnAItIO0PATku6eNPYWPBr3WDp
aWYI5xUcbzSpkxh73VE4POtRvdKPLNtulfZNmXTqQdfpzqDyGfwcdvGJrHookw35HELswJUl5X4Y
9GXnbH1vneCC9uFyf7RvCGr9TugClmJ+MeMDnCPEb2vL1BIM5iBeI7+0rFojJPrYVGvxAuvS+sDg
bcawoBcaNWfDm8+k1neVmqsfaFKIaGvsh5suElnikcnrragUdaYO2wXCXCVPJ1OXa0g8WiB3LGFE
6/n4Npz7IpeH8Ivx5N1GypRSnSXyryk2fnVX/oeKrRnBsisbj+6/scoKlsq95gk3WAeuQjhsbTcu
4AqI06t+h3hkP85rAobiQzjF0gXne24UjPWwSes6ndWxC9rZLqBsDOTj0ydnzipl501VCc5n472q
xUOgCwcKKeVU+1mWExk5DxCJ3tzy6+nX3uUwYAXRoPuBJIU5vm/LSZVtmC7UFx4AbDEOOHDdWoG9
UUaPRPFeKE4m2GwTazAH5zgL7cdY/B1+tDzNhERFrvKf3+RUaPiRcwqrXaeR8MV7C0Y/H6q34fA+
XX45PKLNIZIOpEMZrh2bcZhs+yL0c3VXgQoiSgZkBsR7lbnVdYDXouJNHbRFYW+QILarNDowbIA/
lNAUHKPOdehlicG+nJh/JLISawHkxKxZIX5htJ16SMySE+lkKcsCA6o2qg029+rGdU8CFVlzUWaH
KeQaTOnxhgg5BKxH9OgMtHfd5tlZx/qTj2heZHASWMmsMK5YpZILW9mhDVnbwueFV90sFUZ9vS3A
sEvH7g/EgKat3+n767t6yI6o5h/LxUSd7IqiBUftKiFUge+nbt15mLu9geLabdg0wckZqc9sF0vs
7rQt+V9lbfSXWO1M8nXaxR0DNKZyXVoDQHFb+tITrmVxpwNPMV2CMC8boie/nKxuXIPMUqevKOAf
C3V68ZpJJ48buCBiM3S2djmIBOwxp+vNP34gCoodQaqYnTZibWKYj1wX0tYR6YpduyqkicnLMVfn
05+iv2wqAs0gAhi1mGKLnZSjVe97hNCl9Z6hCEydM9uZqvxg6f88gXWA99C5eSXJCdOx6YtZpuss
AX9z92Nvs1udtGPt36poBCkYqa03CpZIOzj2RHSDkFvEFZaNhT2E5eTV/IZU7wvh/Nou2POo4x7A
PpA+ZbQrk2jdhu4J2vfegMJl39X0IcwZZBwXppExZ13XlIXtZEHRwqhCS788jnxoURyxLxpq4fxz
z97XmD8cDPG+N1FSOxA9nrNnuGeo67+1XhNulYyIxC8WIo4syKfvy80QuYduUAIhejZHKjPKG24H
33goWmT3dtiBXMTylPUW58Pp5BYGCdFfUzwaXCwvjjuMSDitTfkpRK4y5v8/brd9gtsIDRfRYAMp
QeYCIVuEtJ452Fp1WCQiMhRj4tL2aldxZ3tRaKZG1kBFCn9gF6psiLQYbqKMdqeonDxNP5gXxr0s
b841ISDImCftTA2ZxKM/KGbX+vH3hLOEiGDCA/Bt+FpwFGgHkJRdfbmoSSJOWnwx6UpmZvh/+/3/
WgGVpfGiF4Mxjpu4Q9TbzHlZWZlt1NLQmy0U/gyeyPgijavQZVKbNvFO320mnXa1Ya3okGg4JOlR
5FnaDSKUr9IHdz4yqG3xsrwoOdBoI2R+9rAm+yjClGNKSWJWnZ0yw5MWWj7M7cFDs9ie0bgQHRM6
XDSmkWRPWJoOWBNOoMrvm7f1H5I+JoG2AJpNlbfBrohCsHU7jVpvAvgbTJbkbpL2tRKzBi71PrZh
8tUFetjCb+h8u39N1s/GDKa3crNODpMLyachHHEv0KBPucaIgiQypc1u+R/ufbZzQiZISCTMGL0b
wK1qVN1cE5CnV9aK2uhyGvQ+MfuD4d9R7a6wmm+Txv37P1VOVCP1KHWAffqCyHypvVpWzp0XBT7h
HHtK7ETSYOg6f7cCtRjoGkWDPgGrmFQQbALJUepqpUoepsgpoyI51IBrnVDkbeNUNwtEJco1VH0s
oJt2pxbv5XodZMMs6OAxxA7l3SmjEk2cFz/9gK5fr4dLUXn4nSj6dDXBtswN5UkUBWpRZTDDgtXE
cY0ClSof0zMhAXSAc5F6DvFDBQRxY0SQkTrLZ70R9qHPdc5R6wcM0Y0tBd+TLVjRJtmeq/ZmH/Fv
kgKobrsOf/6TiDzaOaB0pP60wD51/VCgP+HSzjZyk6tBqi9lW8Z7bV4CCFZerjj4Sl1G4C1ZmQpu
PCZjf4Zan8gIrrBmQ0HUWbdwc8AXY05m3GnvJjEwiMprI/ZNhTH0gqKwBYwGML1cq3mNUlnKoay+
DqtNYPL2gbjcW6qgB7WPoU4yP0MlKyb8yQZlThN03eMPi58eCFfqq83z6024a/En3Btaq2fEIauq
SMcuCGoF9qdxYURoI8joywxdhcHUD0JCWwABs5PzQlDQ75cljCK/t0U5l0dAoGZdFwOVI1yUhNPY
EKAr6q3pM8zKfLbI8u1ZZyY7bh0jj9+bnVSUFMJlEEuHVBFNt71MnACgWDACatzRQFIOAp3NJPkO
UPvq1alCQK5TW8cBbaVjCafM9nvz7+T/kv98FwMbvjY7RlARGFCV8XnCYyO6J1v6ldQii0xHx34O
W/XXn7uhiJrxz+l1Tka2+UKjkkV7CEYfaXZn5Pwd5D2r3gtfUR3MeBX9g3xQucn1l6NbiQlBsXyR
5wzOjnUSBF6py5yr/QTs8oz3Zm9kspLyK+Jbw/1DGoaCgKI98zaXEOTNnq4Qfi02vFfAnKcsxmgf
zWOIsFk2dhRJ+OQ5oQAwi776LlCk439Oy5gAOQD8SuNdQ71sFqLwTOwseT714A80FTToWRnA1Efs
c4SqBNcVJCFV0ZC/Xlh8eeoHYFCWR5ZFC8BvbkhaOKea0ELt1Z11zQTkPgPWGURHVNxWJgvHc2up
XBHRl9WUWfKHFareWTDAQyHJC/QNJw0IERNudTYCGuR8Z7gGDJslj32jVut9FI8jYarX1vpbMVZA
Fp/ty9g7bApuT/86/MqBTP+qKY/mQ4MTgDaAU87fYD+WhJUUet5Wgqmll96DC7hqFW2qDPBN/bXV
cSCDhyVxa6d0qK/safhwfG/084MsjiyNLPhzrL1NucZWbDlIqJqx/AwiKDv2xOnsqU8PaoF8ZH4C
qrPGoQktjh0mA5DQ482Lvx7+D3xQ8rUdLC9tZzdEwffVuevSFwqsSiz3HBLH1r2xWqerVMQ3CMIl
5TaizlHZXotbUFe5EUpT7nEK6BSUIgAzDggzYf0fS5kahU2vgCv9XnzlxinTS76zqsb3Yb6Da8ur
/9svV/gap5Vl3ig0m8bFSI0n8q1qQFjC9WOzJCme2BTqtb1yCzgYj6OcPNROLg/JsVK+csqnwW0s
MA3u2NM02+oSYMlAuU6ZyqsDU4GCG/ZW0aCc/+9TDVlKVgg8mTvTdpqVtnPjPhvpofpUEJ6xBHfR
KeuGRQsBWLtsHi3SsAostr4/6Au+k6pCkzUF6Bqt9smaq8EiDIEF9cD9L+lzwMCpmicHr2TS3C4b
MFhBgzip5JcvZAM4aRqD+txUJCZXgAUI92A1D2Xnlss1sz/ts/mYJyy9I1wRl4HxkAZDaI+ARWnF
sFhkHJzvMZDgbzCRreggwotaIhrnFZg6kkfUxK/rH9S49K2CFsfeXKR6/hdkEmXy1GjMFuOeOzMw
L+0kp54HaZtdJi0v9ey0tD4bOIq1+ynU7qCQu2OINQVarH6qh4BGvORJTOazW3yqmcXOflKbUk88
h7K/qaVWcQ/Z4FE6HdXMJ9OeLk0B+nMHhdipVVuDcyZIZKItQfMWslQQACbmPnhXs/mSB4CDPjEM
aKy0x7mBXjXCS6v3WJjEm82rll+D6hdSxKITZk2bmJhHeyvRzaBkYoYjJ731Ks7vz9qlfGjzdAx8
PK2qlaX10C2Z9pSW0Ylnb4tO2tBftu2t4DuxZ2Dq5JsuRpMGWGZwmDwam6pV5wx1/tAqUmY6zqty
8xwoss+FHxiKtJFtl/UFNWVNGIo4J446ifkOShL2xjSJuEUnz83Cv8wYetKhoC9EXuzQ/jjI0uE1
XQaKtpPR9pSLttOeC9slTl6QvKXhv0H5kf1E47filvBeZQoreqareim7dm5R4hOm0zLMEKYjxZQb
2kSWuRwk9YlwzIocMeX/NSFyXIpSXh0EohlWZCLI3HpOAoLr55GRbqFEW6JJRrgkdFVauXeOvSNo
9hE+GWo8hMTEi+X5qo2ynwRtGT5N3lkWDyp3DzAl8EqrIRgpKYBhVuIuLL8MLunV4ixt9oUhqvkY
wccGiVDmrv1u7N0vIJMg81qyfBSVWv8RO3KIe54jsxVcR682tqlqHdrkPmdZMrLT2PWNaZQj72jA
WF8onLZSvAKZeNcM5H37O+QaQ0tZC3nO9Trp9htJAIxlznGaZHiy/w7XcolTXc2tflyJf4Q8WomZ
80dSWQgaUQ0xCYqnjkYecuvPCeNWhNtYQxDa7ZhiVgxjau5qMdU297iuyI863f1uCqzdGuy1r05e
HTFUn5KFs6swHgMvphtyJMy6v6t1axYno3xCDxbxi/i/vHfKkrzOUcnGZMKkPKyp628QjIQQ5R9C
1F5yFHXM5IiwtD/VnlachLXEpIDBFvN/8puvs8epycKjLvi6G1zPpole/+dSbrD78TxccfcGBnpO
VygfuhBodFT4yry/9aYY/C8GGztU42Nnuw1VQYUoGLrRnlmeBUjJCoHBW2KxXWFE+d7MX08GWTjf
zuSsb7ESE840WpYCynaS79pRdj9C6PjaJIB4tTpy2luUN0sF+iBGlWco+WDK0imIS+HXcu9QJR1O
dJdIuASOuJ4SEXy1z3C54P4IVVqr0AjcL+wDaUZDELKOcBWLrrbh1kHJ0dFjHghQr1buHf/Y1Gfq
c7lSF95eK0/prbB468m4k28Z0VEYYCl5bt92etqkaxYdIrsRsi53RuWiPd2ql7zf07fKSYFO6Qim
r2ucNv3W68ITRMS/5P0ghjq8OLBtTsqOnKy31UAyNVU8Ck74ke/uCho1J/ubZxrnIFAyJ0hVEtn2
xoV4B8f224CEoHG3NQ+J8pIBDrAyu6CMdiCjQCXTLgyf5QRlY910qyrk62H145LF3x0csKrO/M47
Al6WBZZ76l+o166JEHe6bc1LaeL8ayhkJTaIh5Vz2Uo5ONH0Ze6Tw39eq1brgKdNWcNRu1d5ls8U
UlgW1tvcnl2xdWFyKGI+X6N5gFVfoZSxUqikPxytH1INcE7AcdNcL/lV/j0C0bVBWYoFUZPw/mVE
WJfIbn4LQud3I8wQkmXtTr4fOfaLctN8lxtE/0wjjSKiL2htyw6vS2SIY2rwwYWvCpVSd2y+W3dC
Bsg2G/6xMr4fcO397suN+3YvTFR89pnlaxebDyBVddBLY5mXMl3N8P2pGEdiTET7en6oD/KwYdb3
hszAeW0/my/oB5dbyTW6+Wn0lDcUelQCRMVBPRTFdQjB2KbXRqp4X64hsygWuEXo4Rwx9hpt9+HJ
mBWL3dra0lrERVd6gyBdhAii43Q0XtGpzW9g9zNkz2UFcdcL5/WXLdS4LXw3cmj2bDZhNMiRcpA0
fPku59XbvKCOVQxv8kvDooodXaM8ojpIDgRXF3/Yrcl0mJqb218MBJSrHzel+hBbggT5aWqlCvr8
xchBqmWPiHKIVpSYHlZa9RdrVP8axqk5BgOSWVtDiovP7w20oU4CEpQvkF0aZeqVN7EKD7zDg1NH
ksADasCTuzb5dN58foz5NnBWvE4NA/uzmFPu6UvnkKybqfe2TV4xPs+6x//tpVnsyX1nJR0gQ9s9
9HL2j+50L8dHQxwHHfui5YnA9bLr2YxoIHNZSrBu5cERyG4sZuU3kAgS8RHiEvHAlfPhFkDiDi6j
BDv4N/ViMS2eBKPzVHNa+iJvwKhGL9Bb6MEb4mmJljOoJI4MuUqqLnUq6m130tVp/RlI2ZEg9bKr
0eVl9M3GRN+4GKsWpUn9X0yIKiSUrFsvKYfKrSRViv8okfNp72bgyHC2Ihe9GEOuIQfCMVDubHjJ
zwq+EMi8oDJ6vrRtACi8IrAzbbq9s6dfTsqeQuKBYOtbxYkXBSRQc3ZBhoaB6MEeY+I73V08MJoP
p575BZH78naJPAbeH73wP0/BbnnEr8+FXW/bxwscWa9JNpaIFxr0CkvN5J02vSpO0gtTSnTOhkLY
s8P68199YNdvtAHuZ/HJzAFPoevDFBT658lEPbk9b66Qzq4tR+t2TJcWMKyV8zMmM+aZZTLEnB36
UeSWOc6bedcCOIbOL67n/WT5r/scddF/V0rD09c1vbTPaQjlzn5ozLDfxDvs8q7/E60BEXg5cCAP
3spQwwlQWiDcY5xiOTmkUys4qgSJOoibbwn8U/sEweLGeCq8H91/gEdS0KnJ/tExnnpenNXia0h2
FieAbw/eZlhU5U7J1r+0Qy5xbCT86QvtVlNpd0sTioINrSt/+mQOo9OpV35vZjePy4O6AdBpl2Tb
3iL9JX+IxhEf5OnUVAtvMdX+wC3CnWMmSjF79ZJmT+7pnXaCBYdZQ1hK9yjyApn0bHM0hmO1PQ3q
dC258K8YT0t4Zla082X6y6OLwsi6sketB0ki55P89KzJTgxNhlrbV/EuuKnw+L2+DuKoyFYEWLdl
up+a19pgbS3c1WFM/qcjQf0D3o5BwjvbDWGvHm62VrhbuKrYrkTzDJDDp5LLI1alxj+yf22/LE2F
TOMvdkycsyURS98j7D84AVLwlrAYZf6q/iXGoxiFMZMTm5ocrq1m5Y4PIyQWK0akYNwo8j6J9w/z
CZckc1o6v7FMiIzN0HpKp1Jz/iX/tBmVqutCdrkrYeMdgYDDybipZ6O61HKnZLppkriC0zwBM0p0
7/4QtonvxJRbZZmJlDp5glAdKd+nLrEhs+OTSBric76yVojREXS4uikbCNo3zRm+w8A+q1BylyuN
XpGGj9plwYyZehr86B7NFYwmJPb4Hc+UTdMbxjq5x88V2+tVS3+mW5NMF4dU8UZfKEuQqBHPZaC0
BpmpdYZ6uo7UdKBQCtofasBeRfgJsU51VRuufZStkwal8hLNvvSda30QXkqoUFRHEMVMoJKalfQS
5BOizNKkyYib0AgVUXgeOIRq+qunY+rJWOn4P1IZPHXyUppOxjCi0XsbOfiazQlUylAsibqJfbIl
WuK/nV4YasFBNVDfizqM0AVkkTOUJ5m+9iNKX2u/LN9LcOIPJ5ukFl7hhRNyXFbiioHw+RY1Yeus
brzRaKhk0qW7jSbDju9EjIOiV+vLnsFOgbmbenAi+cc07O6ySgc/ui7WC3DrDPMWYdafKfOmVPRN
PrSpk6xETd+sSa3MAvNj7vp98yDzsbbGW1qC0KNybTMvfVxxcqafu9HaQuO1ieOBDtkNnffpjH9T
5Z69k0dUe9Gcf2JoiZyB7kI1DGT+E9j8G3U5hF4jjjefbSZcAu6Xg3PODdRTQUFZhp859W59acoC
xImWJId/WCsyGMrBG77HBIwA7/4SW4avdHD9J3P61EutL3rvzszSamtIgemw3p4DdH+dTp5JtjiA
51XXhce45R38nBk9VGE6ojYclqBNfO4S6R2VJIPjEnL3s4RgQj9w81ShZ38YP0cVhmk0oDoPcmOL
DcUXBgTQL++IFp61iG9U2RO+I95B46n2aPF8IjXgAiVIOvL/nWy4QaupdVB0I2nMm57CKWB8+qfj
WqXbRCwTRVOQutDn/dFp02f9w9bV9y8dy9bATggxHda85MdGAjwV4MLBZXPNWwzw3x6zBJV0teOX
qqYHPryUtP1Ey6GJQ2JcC335OIC1A72GM9sCWZZWE0Atheu2rICJuvRJQCZm6I/DvKeohrx0n+Lz
lQxkciIm8mZsmcjNFzI976Yj95Jy5OOCklBM3oJaq2IJ7g6lFakTX2xnzj49peXtrhVqsHT379qa
NwU7Pr77lTN0WfOq7t9uAmzAc+CLLuOPYbpvv042B0BQHxFgRGXj7ArgC//qIrgcUV1+wzXVHQVD
OpfGIBPfHxrKNgVOK5WV/qU+n2JEjkHPeXCulJG9s8BhZSEFXL5dM0udO4HjMA+U0xubrI8MC8Od
y/qUzniZLl6HNVhWa82myc/gbM9UUQD3AcKL68nxnObp/UMy2VnmZ5VdZRrZ0vsKPJjIWEsHrj4Q
PKr1y4onPMGhKGypDyeeOSJz6bCrSuAUfdmnraRtv2hwHQNah4n+4ihg1Pz3CpM0rc24OPPFCzZc
AHqZv47cUYoTbnQmrFXiZaMNUbzPXcj9BcI1wBV7TFprcqA6lGNiNpw9U6sYc6L7j3bsXWdHa/1J
cEhoYUwAGRYN0lbv+dt+FtJ2SXnh8Nv9sltTvkovjYuUNVRZMrz0EUqdsc7dPGueE1wsr7/BT9np
GdJg9uN3/gCRfsEQYWoWekqJynp+3jhQPAhq2eta+adUj5J8b8h34Yo9yW5h08c4hBsHe+EqkpX8
BOPXEjdj4Cq7QTsNaKgS6mqd2DQlREKfWgQOHTHq+rxa09W+vTMm55TMnsVYE2NRUpL80Q2FqIUD
7gsXNETlILUsm8J5WCbgZ34Gd66JGnkB4S/nfSzqfrDMX3Y19pA3FfxF9YK2EQ+dxyg1mryWqygd
RtO8AJAf9hZih5n5ft7uyS3weWjv2AGW6Ojm+8XkdNcuQG1uaBNmhu17LBzJLmZufAzKxM1UNdnD
aYiAv44ZsDreynax2ZjDWfk7tkp7cYPxkdJJS87WApKBNwOe4I4I5Nab7D3P5EFyuMTZ3oKuDJ4a
cW6+Ngl/F/0kZd1GCGLpt6LD7yfWnrhoZem8rqqcdin411rDhzhXLTvI00AT6vCNvXDmPFNF+Iq0
NdEG3BEdZU6Ov5a0+VpcTeztFS9gZWoCJSeQ5gmU0JXslZ1RaeQHwNKRhSBi0I1rY+JJFZ9aK9uj
IBsfVen9ODQRSC/LnPruWxIJmbN5dS3u+U4L3Ik74ZKrgnUoPf+vTDU/qttx/uRGcPEZs0KeKhYh
Q5BbofcgW+i/Q40R0ZPOa4wYWLmhIdDFpb4A3VLGKiNqkY6dutbJf9xIDxo7jd2K8OiI4GH/MeRz
Q8gwtLQNuhGknV1ba96sSfN7ZYJ2JApP/5Nw04YzgHrNBysJRbWO8Q88sEosgjdXf+hxN/P4XBr/
CKXRNJ8SCzrFS37dndsNeg4kmkXLtx7OXkgdvcOqwSU7mBHUSLZr/t6fvkH33JKNVxzS/ZaL5YOU
ypLl1Gzsq5eJvlaMhX8GH9J6c/u0c/NkXDX7lAknROW7KiDbqvoNk5SkjM/n6bOC+LtXtHF7y6El
TjdBFOWOvKIqvCqSbHabX3oBeDcJxvqhP/bhPhw7DuHO3pywU2D2GFgexNF02RoGgeonKjimfA8n
ATkI9sNAB32Tgws4tVqUFfcCy7jPUST4NK7VJY8N8tKhuhmkitMaIOY/uz2MYFDDRUvbFeOASkdx
7l4jaNoSjjIqZ483m+pZ+w6ouirxynzVpCkmLLY0+izH8PcCTEwqN6Ku9Y/6Yup473IESfQmj+dj
1idWOzWW1iD6TN2122uChen10EwNQIYVzuEMsV9kGhyqadHarvDQlUBFNDyX0eQe0ZM0jk+pk1yV
T89daCISwCVnKAjNs+Ydxao2YUCr5nd0eBt2DFmp9sMR5VlgUEA6uC/uZOiB414mdaJR/KIeDwW/
mH5m3LEdndtRqMTT31g4Y0kNhxpVDYNNdcAQeBHDNBVgaWkyPWzRZciroAJdUkXqjf0YrOfXncRw
7Z0CJLoSQwxqjPe0nE9o8pKH3Py3HRj768ueGIhGLi3Q3nkIjxYoEeHvmG3+RWcqwBx7phEwjWoa
Dx0Trnk9ubR7pheFqwrs/zjQiC7p6cgom3hv5yhtFxyUG7SLOLodxbGQtOp9HtweO2cCGC/yR5A0
50dRB8z0kOy8vzCAQw3eo37Dneth8lQNVV8GxvGqhYrm9V8swSyOdrz5DArtb8Re1MgRTtDW/rsL
ql6TKAiqUaC9osjAgpeUqf4RUuWVrdaPzyFabh/8/Wne3IfJ8OIpBA0ywoZd60Xsazp91XtQrego
fATwo2/ko4WXu8ZIf1wVo9KODOJ9XuJuWEaGvKaodYNRq3tZTlZe375ubo8GxzwOqPYTaNQmfBxQ
aUYti1bU0V6J6FPJxFDtzNfxRVsGVt2ISbgyJoHe5cw1CfNfhsL8jDkiJWERNEejUI41NFU49k2Q
YQeDAbMkZ7xhRl716pDvb35+OQFZ/PrAnV3MJN9Wh3mMGTATDQZisloje6JVZ1WD62/PX2Tbam+R
MC0srlEQpg7z6Re4VXPQb+m5zDvaiaZAFFsWkotKe+qOg/nU/9VVVHx4Oj/ZPC8u/cbQ9sz9AgEB
31kI/+Y15dgMmOl72DiHC8LZgLNLoMxVCOTs01jYPj5YIy/44/bnYJtHWJLIl/8/AN179CN34ZL/
ShF2Wau1hS+w7w8CreRky+gVn2DbRNSsVnhQrnqrwNWLBGDda3sDNJtDAiN+5D/go7NFBwlBsKTT
+t5JkT1DiHis5oIjLr0Ol0lA/5431SOynhIH1aPT3AkM8tsN7MFqOyshvfuaH/AalnbtuE4UzpJZ
WLVOx1RmNUcWx84f4XFtDw25a2ICVlS+jSPU68bN9Zsudz8PChO0TKZWpenDZT/oKPW+KK+q7DtS
wWvAcBVEUFcyC3O3TgyZXPJRrYZWOZ7Nw3X2A6uG3wqWVFH6ROrYdl5uOi6sHl53IGwSjZqYsS83
0Hg0CosFL6E0s7x/qCTfnYeXLYzc5MEd6dGqP8T0uGX9YiurncT6vIWVeym1xDMOjCFMxjHvoSED
+Bio4zGqHa9eqIL6bAkCDJJYR3JKb5JYhxTWCONavlb83BSvQgzAmHkyqOMHgSWbGkSu8qtF7kix
40Scb+taPEPVe5Idd0lEYnP1PIoZUxK2c3NiGc/qGany69jQzeDHOcz2fqNbjIHEDOrqYtRnqKT2
iQk2fC5/S6ft7IE2YHinTR05GwNxi8XCl0IOMW7OFwMmJDEwJehHLDDPFmQALIrULcvEP7FAJr7U
58zBGQstf9+DzcUDu/bq2Kj8M7MusVTy98lwQfzKyiBde9PIVApJIeF3M+FtdVyaNIkdGQOYDQX8
q5e8q6jBFVXkM234PzuniwDwZpEvfjo5iovLZjg2O3WfM98ZC2CCT7KjonscbsOxPnB3A4z9AqOL
jsDMKZpwBnTjeh+pn3sgZVjeZPkXMd9nnIyaeu87nG5XM/ud7Rz49aZhUdTMQ3+I/4HV+zDUWHcO
dQEwL6ApppYufrbbdCr/YUJd017S2Nvk7YBNzgro9gHp01DEAuwQoq6z4vks7xwp0qI8Hw4hjM8z
MFPqijvtJqZNAD8BxvXcJ/GWNzCeoBpQjjMGXGznEwcIJjynqfbA0UN2qaiet34W9jC111IgSXIX
MKjWU3M8W+KAItbbuS2ey1OlU3VVRzdZqnkD5rTSXDedukB87P6GjAZkPMQeE/3bcygAph0SPQVw
ntzRnm0xSOM4jelzfc7kqyl3QObYEiloxc2UVgHX8b+2HQ8sg8wBqG+W8btw3ZJQ3i7YML4eKAIt
wbm/0bccBcCqCIEUUD/Ik1v8pNCedBE1wHOBkI+GKudeBH2GGocjRglPpBCTFbCJb8h/apJ/rh7r
sggmm+SrR3kvDDhmzWFiMw+aQHQLHI9SC6GDvjqvJCw55OCOlYmqNP7l33f+RcbZykEqboHpHEtd
eFPFFe8nAfr+5Yw9igG+bLEhTOrTxprfhIHRPjQLJOnkU308irYvj70lpPpjKYiatL1XCXRcNRhh
wOw2MBlKynuJlPRPUx0C0uph5Ga7kTUAAqh3y6FCM5IAVHbGvisWQJEcsLDmk80wUHxjIxuKv5o6
d419JNFhhWqRwOqctpM/Ex7DdwTPauKmSYklAe4Ex5BwuTz9Azv3pFliVIemQ3tJGzbUtI6bLcLx
DAekPg7wgogecbrm3nJcdsSEWZ3tovb5yLI/RuUu8OIRdt0W6wZibciIoDSxsfMmJ8djxni39dho
FojkXNqrK+Cwy1psUFvc+UXUcW9nxHAoSOmT/3wuWot8kqMoIjw3aewuR1J82rd3XzQ1/kJtWQVb
twGU5nL4p7n+A4jVdeTS4dkN/+W8DXk9BsH2LjLp69FlylZC0v8bvf+PGw2K4XPokETCP3gIxeZk
cllyyFR669z1V++tNH63SgSinO4rpr9aN3ZY3yT7L1AkGtcFzl1MoOyYvHRMWPMpxO9MYM70ZgIi
ymNahqylVXIOWN56u4XCTKfpIOY2zjI6384FKUWsE2yGtDlQFZNZQvR/VljH2tckHPvkGZhRPYC2
2cbl0X9fq4SDTStRT+rZ7/aVdkUOS97bQ+kga23GT53LgL0SKLhHXqO828Mb8DAlNtWTX+o9yKj/
/YCBqoiK0ey8M7Yze7cINSvaPkIc44jzKMDjatlvyQlRtLEYYFsTdiQYdREa8ZlZiXwkbBo0EqkU
WUCtZXL7NSqGoSkGFT6fePKUQSktsvFlDVN/CTFBe4DuqTtdLBFnM2ZKh4r++92YS0VE0Gg/Oyv7
XxPCtq8iPfDQ1NV6Kyor/9fYR6PFynY63wJFYcfJXmQhz6KvetOdQQb7Qs/z+Fa5dchjBos0yX8+
N3hDpdmmmdurhJUB4tIi46bdysCstFqaN1Mwn9lqgvsGr65ed+7YlnyH7HMp/QiUcXLOPMu6OxR6
/i0wocJ12dL1K5kkle9VqxT0LzlHy/QsxQUOXzsoVazT9MNeEky5sGiVRDW17blnQ/q0gqhDDZJ5
4nnPsBnNn6kgGSMVjOiS72vLNMl1y20Z1O/0XN89ZrQa9XIW0uAmE6XYRFX65rayUmP7lqjUkoKW
FOChgoVmAzCnDL0aeyuPZsT9bqooXNvboqN4Vfd2gJxckUGNNUUl7YbqDABJdd1a2s+KTO4Qe/7/
oVZCq3lT/Kv8Ks6MSwvf9dovziQ4T4kSrfhwsTO5p8xUp56QUTeCkqKJmIuoNLYVZAKVtWwqesqg
TKGSS9wrsesvcKSZ4zr58RDWUEo1lSfA25HQe1GdL8vw0bsZMMpaKy8Ld31MW6I0zYj9h60pIIey
ph+qoday+yguX8RoJPKfAq6ElMqx7j8Gkg3b5rBVIPsNwp7azXVTY0oc/LSzF+gVldCKb1SiaY3o
4xlc2EcZhr+a9TjBopMgy0cSkDxZFi04D747i75G9CUpCZyx0vVGEKjTtuAoJ2Ye5aUwSnH1PYRB
mxe1ryp2y2GHfI5vTqI4OqKyVVkDxsItkuCRlIAX314gAv12eNTs5rggqNzhzP6O15s+llmTONWq
N0C+U7ia/Oy4hAtJSrt7pV0VZQx60caK5p/lI8xHOOKeVPaPxnNsRVtHCsAemKBDKUmcJ6dzOn/m
gDRn4C7n7CD2+tM3o2UWmZyOXO5Wn0SvZj77990F4LP2kopSo3TJfDMsK9K4tUMKcJU3dHMr8udZ
bVX7pTmH5nI7TivUCP3GJALglTNPOFgjg4r5KPm1w8zK4SVnUlVtgCxeE1rWrckw8OQUp+VFpuDc
7/F0ihfOHiKdign5DR/9EibdXf6TfgFjr8/dmzLAwSvDLx2GP7g8M13HR1h6Ti1uZ47Es5s8MMsI
GMYusXLshW5qV7LQaAkohgVcjaGPlO8mMC2JTFpmK5B1Sb2TPOZUz3KR/LXcvV/eWF5BdsCTMmg4
LuBI/qAjKsJaHtAbHZfSHazVW787o//g7VODVuMCG9t1KdwgzsF0Rz1wU1CaleW7wJqz++rnQFAE
3UegAwlTgUTqZo5Jc7Kua9+dZGKyQIh4pQX0WHmqIn3fiVDlZVJRIZzVbb/jvHgr4cMZ/luTmN/c
1q5RyF/sdVkFH+UKeiES1FzRkqujyE6MbRH1L1jwm5UU7a514tA0GMe0UYegwimjbKftfvgWlZ9v
jneSlBHYfDxZI6xBbL5kTqakzG2SeHh9XVvvib2WcT7C28oleeJHVGU5Gm6VqZ+1UoL2hn7nDAXz
CQgvWtF0sjYrA0w1iMOttJRg7lPdzDsKW7OjMj4wUE9q6PwOWsTabUeWeuwrcd53H5HJJHtrt7sb
JK51BdTDRAqjtmVZhB151/e0yoWPWOXALwqXuhhSBARh0rlcbyLFk1FxfglH1nrK7vOYnb91ODPt
j17oXc9y3yzXtfro+k8szyhmQooMCmyW+UdQaJZYn+60E8QRszyAj2s2Cfz99zzVXxcREUq4H6tJ
c8d/Ymwyl/3fggyDYFpon0Fa3NY5VYOnIW53dC79xn5TqVjqcETJSiM52SuPJsczWQw8MsTp0oPt
A0Biigtb9MUo+wxtp4NkEYrBFeFrGb8NowOjjrFu9BmxsvISmxLV+JZ/ony6k28iv1fj4m5WMOos
Cw/K/k94m1ukRocq5ZxDLhCHz8yC2OJvc+gkQVUmt85QwTezAAHyWC1D6eOWJv9QrA4ZXB9jOniz
BCWav9b9lAlx7yMH+DXsrrLkd3tmaB2vB2NwW87Zc7sVts8cLWWTASJ2biQmsKDAK2yaH/8qzefi
0WKTkcNa5rTcVxiRhHbdVuEITatKQ3QRE+0ByE5ay1WTPf9C2MO0urXBE+JWrqwi/P7T6/MvGpAG
GBkDvnPYi97leCIN4uKWGtR8uMcPSEhSQTK5rh146WseFSQt7BSE2Ej7vcM+BU23XQ/ZVk4SoZb0
DSUAfJDAtCawJkTKfxEpzQtlEpKgd646uE56PSpNMRjm64E/i0CCWN3b/DxBwlCO2j5Ve4XBmcLo
PineuUCuvrXz98YMit+AXR2bWTtMK6CJ4/+jWHUA1+JqL5Tzbl+Ekji0Ww3rrn7tCCfBctMHTuiH
dn3SLSoXy3bcrLIr/YE57wUIIy0L/+rda7Hg0SFz/cBewhmwKpE/KA96T1jX0VJmzUPTMC9OfzCe
/ZMOFLBtSn6uYbhKYqPmQ+TbBfrtWTF1MJiv+SLbPtpfF4NqiGtlndGSpE5qKm5vh8UbKDNXncgU
PjjB1ier0jDr994xCtOFwhRUEnGPLc47yohDfU4OO/aqkUIbGHjIMPvpmR/eEtsokhAfmKIETcOi
C0/32rQNtfzV7SWPOyhXvi9YZyEt4Lecwu8iwWaV9hsgO0zdGSpyfFz17uP4MtnNkCSo/KOgu2v4
u2vn1wgM8GKegzJtiEXvwIT773+Xb4PXv2JgoqwtqTASyicMM3677yE8nSa8cE1H7+R8PkK2rQHc
mDzpAPQoj196fGV3lFjjzXUiDxczNqQYSRaPg4uqog9XkjpvsnpgTThgTYD0UJl5DzwUdkjsK0v3
63kPeY+EfDUKqKQnqiEdNiEmyvrSnQ4Dy6LEZBEUW4QlcRK7hFXb/D97q6ys8EGJUF1UeTxlI5zQ
+AjtsrA9BZ2w92IxeOzR+UO0/cAMuPbVNSY2AN9/KRwjv4RdvxKLyhYVsuR8laR5qz3vlCYVrEMJ
cu8+/FKom9JNMrbDWcwQKa5BgL2Xs/ePHC+0RRgWEmpn7tdWUvEwJpy6i07r5ZwyA5xqj78UX6qZ
CG+h0EfDR/oyTZ1t07TZAmWztq4lHArMS3uRhgHQz6d4vPDn1vXyHtE0H5aHRxmqu384Mqgr2nRN
ivfI2h2rz8xjAzvz5vqGdDWFXtCJe70AIBwNbrxayKouEOIViBLwi6CvqKvuvKUDUyIG7M2bO20Y
Uv68JFtzv2dQeYkrEBnGbU9ef0OgPRAIlPueB9+iQegBIpjqq6I9sV/HY5W35yXq0lOE/YQDmz03
vu/bXg0eY0KCB3Vvx/ca13SzsxzicytlPQLSXXqSwzpuKCb4bAO5JuTX0Eq+s5VqOw/IgJOKzs1m
2rRr4AWzocCpavIllD2xOZFVczofDSjzyZAP7X0j8+PLUqUleaA+Wu8sgArR9c9jUoUenYO5AEbh
BRjunu04xpES/VLTa1w7NzaZ6kO9oLkOHusCmTwL+tjiolMQWIBce5FrXaoxxVNG1udYd0djIZZ5
/e8fg/ZnDSWmlgLHyxdAMvEe5ttOFFuuzcq6F7Jv3bhJwQzHGoTmnU2/qFOjFxaBndyq5IbPdAZ/
sfm+hyF9xLOqnqiCLPmY56XMgYepON4PoYu0N0l6/7tRY1hr9LtnHPM6pD2p3c+hgv9sJZWCHnOq
bWDivK03eCT8Vqx3ZRNWiuzLQak9gqg4G2TBe0qaiWMRbZPAxLsM5AznYHTGzAQuVr+npAl2xdbz
zqAVbqbaJame5bIv1FMw5FeY9An2X/RKo6GXlnix9mipuYa5J6Gl1f6KBglPV3n51ARKAeP/S29W
1YWAKWXVbUnNttOpTTAS6CVqJztyFSIhmlP2L5+i3uCebfctZQhOuEBei6JakEKdqpq3tu/er/4S
yy4KG9tyrrERftfIvatw6BVCQxl0Q1SnR7hIAgxK13pNWQ288gGeqGfIMAIItvdFNOk5w/H31qJ8
x48gbBpI3KHF3bktDdmcBvzxjVPgzKS5mmfZbT5ZK/bloEGr2/1uTOWLoCs/+kgt92R+1LbJXCT/
CDV/FoyiowWFlL+x0TV2hDf9Qe/Er95uIOve/vg/aabkWCrzEBU0bBa6bxKK8hCmazZ+Khp6/vmf
HkvpSjPQhbrNbJfLPHG1GyuMZwwLGC614D0NFay9QrzZTcBJqAaSxM1MWbhxvBHLtAgWgJYEpz9S
dzqJ4Yl7QdCXoOWnFFUp1Wrdp919A+Owv261H6lt4oaneoTDzUWHmyR2A7STnZnnpuObL07Znfty
sfR79H9tTVEsv7wMWeqVADYCnBHUv0BhseXgh2+HMTY0Pri2Bc509nd88rSsVXqB9e0pXyi2wOYr
t+mpei8Q5HCuFmWLDHt33xarmyDqusrjgteDxs12LhVQj9QmBiuHocIYSbD3Ss3nOZYEz0nsU3IL
/SmNRHN/CQ9ZT5nwnL4roiMePON7WFuxnoBQk8B5cX++uw3e+xekEWdu5K4nwac31/U2AFaiAb/b
QQZqwAFCd3sxL2mTYRUqVNgxQUA55DzAnuLa6OFC8vkQUif7eKBDuQgAC2CgAFS7lJZXOexC0ffr
mKueuBNNzrF0AXqUHTBvmBh3wnCPATGEnD5tR05NUEmUxN5aa0ADtRWJ5OlX5Ss3iu7DlDZrOAbE
kqn97i5MGbYahHTAh8RJIyY/3vWE2CKqmdRW9rLc3kcP9QncBubjw1L0i6iFnvB3PEExoGZVNtlb
2ao4QrdOyxwXy+2f+3YnzsM2p5bIECtEvXX7yCkTgNMSS5WJQk40PgH4FBwh8LNSZl0huduAN4Js
7zCtdz07hgb4lZH+KY9XbJJSP87TurLqQ3immo8LgyvkSXSVFDAAp7DDEQP2CjEYVO4F1/NlVruE
JxCv08I97vwnuXHvB7X4pzwo3jqgrhwCiBlYTRz+YH67SgtGAopJHW60QWjFFOmaStLeeNBfN+fX
07yJpFisU78BIedZa76q0bbS/UtOcwDoAyEm4zJqbQ2lu/pvUQqNg/ObmIgUsVEAyunmID8I1KCK
JZpGqHH59q8LyfROg34wj5ISlMPZkXYwKximcGQH0oROCUnPHmd13knpX1cp9QoSOcyYHy+wujmB
YxvQYHUVoi47YXv8dqEDkHgLcr/X/nx0eEg3mT0EvQ3iOX345b4krOfS9txwy4N9iVnWBOWr5VWw
Mv5JtxABXPm2GBzhfkjrYC4pUuD2Ptdw+7mb81L3ava4LTWUYLo1/d026AKN+OqwAs+bcBWMsVUJ
bec44ZIV36L5gVO5C2SKql7IDx3iG0z3259Mb/sPh1FpmDpFy8pNwELnS+mdWATqz6LnFsUrcozm
sItFZTh9a67TpbLqK1m0WNSEfj9Yt06USMY1FqcoBFrfIqjjIB8XJIAURczQHKNc1QyfD8P1iBZ1
m4F+JGVLbDsBje40Q5KNj/DrS1ynCvAxc71RhOvGN4skmFwH5cJkfk/Sv0E/P7zbLqk4/UB515yd
f0jDrOJIbdv3/VP9Xd7my/SAh6G1UlnPyRiyGDhj/Q1qim8LNm4E6yhPnDh+bz/BvbQC1uG3FaFs
/M+6sajMn3cK+iUm6cTfv4ySVeG1ZcYylpTlIlsx50nJL5q2tShm9EYSMK7ZefDI/uwZtBhOEsPQ
pPXpeGNEjxTpa6Xy8VNHU9qlX5Qka9eJq4wARAvhKUQFAANh4Kxs+okXTfAaXMYyImJ8Gy9OIkBC
Jv2tJv8im318F1N7ZbfN29L+bLj9YWWjtD8eBypjAUlo6qAUx4Ie96+sRHl9kulANS2G9OnkDd22
EIzXU2n6UAbsN7Ety3cWwSkuOmHDegOhW1I4DE9GVBjC+L8l6/G6wA+ooIbsV/oRMS9vp4wDgsXt
bLfDMLzpIfR/FpdtTzTK1rjbKVB5CBl4yQjXYpyulqECmPxuOTPFer8JJNkUq47sIny4IKQs++Ru
Ct+mbmysd1+v64oM7tk6+/pNJrdGygk2sbqZYhZkmlWeW7G5qCdDiSqiPPzB5aibjFbXQQqk/m2g
eZKLEb5EV8dvUnnKguGZp2H4G6hH6yD3QfVHHHOi3N0481LLxvX88vr4yq2gIod1yiPQCI0yM/NV
mZFJqZWpel3JUzYut5GF5vrMXCD4fYP6Zdtx5PEewqMX5qkuMbSRkwnkedKFvTxACOvN6f8VIcLQ
WTJ7WRffrRNS/tpZ/jknNBvQsDREazQ/oEgzXT4/05+ulgFV2ucpya0R/bUHAazJ6Tyj/Tk/Boep
arjoVOvZuc6KY8FerO4kUwq67zkFzJ6yzu99X7/cEM7BFaED1PmQ7/HQ+9bWDx7hCgtTR+vbCx+e
g5ZR6bdPaHC8OOg1g6yT+AIT1L9pMOwOx73v5HGqyUjvtjGnfKq1OiiFR2+fjehmRcggMHTG72AH
tvO7aJi7Ink31rff3ycOrT6zYhX6diAd/hetQ4Jj4gd2xcrj4lH5anoi8Bf+hu4zvIiDnKLIXQFl
WLB/GiEisoRpggCH7V8XubLFPA+FACLIvq+8ymXSRv5LNHwE5aAfZ7AEtyIhsJftDTd3Ng2xonEI
QHJtOSCxzliQpvEAYBWFBgyuiWs0Rjn2UXmUFXrR4KBRszFcIX0JH8y/tANWwLjPb0vcmmlf2P4b
64jz3vVG+Daeo9fSBLjcB6lgezn/tKxJGmqGv3YqqlTANZ004SL0JEyj3DMPSjvDtLbKPWe58jqf
PUIhQB1Mahh2ILY4EPDxO561mEfMNBnTNHuztZ4QzjFreyVf0HGLBRLoAIC0LLt8h0Mc7VjesVw7
V9oAz6zxAYfb3m+1AXX+khF/U8E4dR2EIhToUY1fQDIm417wF5BgGWfMwVYd1MtYh3jYXnUaIGTZ
kpRLL4QGgx/yfH/QUsOVKjEMPmQSNrIw8gbpPqc2Oi4sObDBZUN1GFcpeIH65OsqyqctZsowUYSC
jpRg0OXVhLLXRG+UzjUR6RTWVsuhT2hYYs6bdxEKJjLr6QjTLFDc0fMywA8OI7msLUzHlg+BcJlx
XHdR/rdc0ii5dZsD/o4pdo0dUkBmaEyX//Mo9VRwfsOVS6Km0AszinDXwNaRCTfHxFLPOhhZofkc
y6kbuOuzLhJ3tTGtPHoC+1Ru2U2rPk5VhKw+M066OqtriTeUGH6G9xtMRFeefAt0wmKqEzGo/8dw
VgfaKZwDKe7NJvTuduPnR9Y2hVYFeU/UK6TiJN8x9XO3VNhG4ijEMvOWzv3tQfs46LJXq1zRkCd8
OhjYCrSDq597eG8PQDevywkZVkYvY0ojDTJZS44KBkprrwBaqhjkJbcnH7foGr/pXeBrgPDCpYX3
CJ4go5e9IHs1WsU7fhfdlQWBwH0hH6KGGwpsw0+D0i2Hf2fw8RcKvC6+YoU406iWm+ByBc47C8bR
SBzYkkIMfzrAZQwoU4hqtF5o2xINHd6HSblw0SSQ2rT/AOYVl8wK0zepEgezd/Pj0CuIqN1KZYqY
610N5F0uGuw/i7WZCkmm/kOJYeI/CKimyJg4h1G2H259k4Am+WDsFA70q9W9J05s6r7poNfF2xhz
6k1ro/hREvSL8eKDpRAEj7xZMPq3/JUhJmEqJP3vxQmdN43DUlUghqOcUP8mjE316I+SkkohLOXC
XW6vF3adWRM4vTLoK4n+uyDvVGa2ffWlHyg/y0Ud95+0VA/XDu4dPxv8CNZWCpx9uOSvoAD2GwAn
VCGroQXz/NSQo4/z4U7/wS+A8gPVTb0RHbFKQsF3dZe3lzI6qdaCN3WQmn5XeD8LDz4EbCmhK36E
sxqz6IgPduAqOi8umB4lPVZHk+GQwxuSoKKHShAIFNTTUyURxdivTKJFdEsT3cxcC5kJeBPEv/HT
7x4GDFgd9v3ho6iA14wi8oCRsAPloY2UTo2QSacDt3dt0lu5OMXTNjlo6YfWcyywhvdZtxSOkHUp
ylRpOaIttBfJjZIplZ+Eqa+KRm+MgslBmm6sut5vEuW2hYK2BDHiYx1S2pMAUCLQLLU0MjVQkzi/
lqhzeFfVwIVRCrgvGR461nRmxJWsb/ORZqowKChSSi3yZzluz7I4TCUUKQ1Owpkxln2Yu7YWn4cl
uXZogk6uAwJfkoUWy2kDXn2OkufxZlTWsmiT0iNOZFuMU5FDXRJsVLWeNXESy7RQy44wp58KGkT3
0Exl3NWPKj/BTVgUarjbEdVb02+mJ9PKmjRr8GQc4MbduWu0oC40YeOj2ybwqxp5P7RK2naundxe
8srO+r2JgevXXrVbF5c4XfDdon6mJYfvVs4NYsqfC2NPJqGGYe3nMSd2RMyyPfcHxYkRkI9BCNHP
bDX6eA44/eWZBR16EcQ1toi5ejVCw6jFavcvbxRvB7SqPpJlm/yY2Ga83O4SVpwsLUHS87t50o2o
BnINTES57vBVsR2ZS6gJWn08Bdj3lVrYrhhgfWlurX/Uc++iSny/mCH/u7f/BG0N4Scqc6oSyyu2
Ll3o/j1+b0GOVlJcuntl4RdDBKz8bQ89ZfSaMXyRvK+DgBo4WJAxdWzrgXP8zvm++Q9HPZgGnUN2
6dMdgCrUqpH2RX8XbyPq8rShKTd5Bt3VHrF6Szgs32CvIYXcz19zkvWiS5RRbi9DQA0y9xl+1m+e
19v7C7Fc/k9bCyoaiDOQ6w1B/3pBlEX1VD1zgiV7kPn8PsT1e2IHsocPL9GadHeLDVXqHtDTvGAc
M5BwKycyfHQGMqgkbylyAYZTX4MNPqICUeDZ/R69tPS9MlNIaUAvWp8HnxitmGDi44IHAvpCMJ4d
NumQcwTLf5PTs6wjCZ4+GlCauTZLOmDUB7+qrnDm1MtnMwX0g3HOS4kTIg/V7bi8LMXRzOQFB6KX
BW+ZcHnjYEMK/koeI6VKa+NFX/m+jFNFXF3CNv7qmBjk1wcxG/j23Rt1BhNLTpRCErCz+miCFTaF
uQMir41SbwjaqiLuIu3jyBDHXwtrr+XAYRfqY/5Q4pPNQTkkMwyb0XcT/D1U/5xnyYLW3wYwgTRk
N99RgGGq6/41TLW2z708NpS5hk7QsOZ+yIjHkRz4F4yWHYaYlCPYZCLKxLINm4Uq7sJvyVvZV2/K
zqoiScTJpmD3uPJ7gR8do11VSrSh8Oq7endZ73/m2xRn5Facs5Z5IdxE5/G8bVpIHnN/X0l16rKC
P09g9zIN0G+v2IEDzmnwI6jMW5aTpmEJNOuzQQE1gnw+TeN/tNPKN277yDGt10HZ8IGbJA0BsSPD
0yihKy/ZaFWudmJ9/fktkWqHSzUj7dppPgo6jNmBN1bHxT5ErNeEpFxqCTBgrMxrwcACKf7cWJWc
Y2u92lidysrFk0edireYJEtPy23Ptw7KZAnr/CN7UCeZ5E0xZKnFsXWtkH5vz7hs2sCf0Zio/Tt7
nGXgjJgOj2AlSlJFmq621I/pGviYx4jWavoZsq5iONpgiT8sjsfCieBG5jKtF5QS8ufSqLhEFNmH
/0KQnB9YvtdL8PnEQI1eJlyagD0dvxfgauEKQyDcOHFHfeNdjBa+3ZDqINq9CH/min7ErdemLXoR
njtac/kSAbQ7QlVYTXfFUKG8Y8hCNTe10fhcAxw/Mh3zRrQpfuWUTXwiLLK2bo0fUNMdpRo2qFjv
s9ftVpKsBHEp06p9Bu9Tt3KnWRv13HiVpwWSc0Jf/ISakbXIFNu0ZNQ4Ice8tZoUyI+SMN2unhF6
UXI7RFN9y/OAQM/jceLh8ADZ4NMeQWBd/ldtzso827Dgxt0g9hvLLDOgbQ+qETPH+ZAsY88ydihf
36SGxOVHLSGYwNUggFZawWLG1uJCpAl+5gRSSS1Wc4/LIO+7a+9q49PBLAW7fuvopSF37TgBcIGd
pdlbfVzOtDqanGdcDHb9hrbQtBvlQbnYm1jlfuLC0j5KsUgqfdISRxsvDSATRS6h7MRi3YBNDTSS
gpX1EwobNf/uE5PU85S1ZwspEkmZt6JgQG8QosCGpWYxiYyJWux0WbVUGcjbjStOVy4FZI/B2SA7
3DAP2Nydfh4AC6N/Nu5cQWRTvltuIer5t626mgQXabZqnX8qHrXlqRKbn1udzbtgUD+0UJbohc9c
8uvYV4kZqpE6olZjkjbuWCTp5uZRdUJNkXdGH28sZIrW3PmQcwJtdaP7UBBsU+eXv1xq4TELIRkT
odfyvPGPXtk3s6nTHG7OHpfXeScMUpVklBzS6S4tnVChjRKyfzqBP3/KZEM23MoAehEK/DZWGYlu
bpXumko6EnHzvsmkZXyMqatG/dDPrNEGfTJTxiQ2QODY0zyCUMOkzrKTT4lYVfZfEdqPo5XLHBSB
emnSE2dTi9B5pKm+q6dh5FsnIW2s9FnvhjW7e0/uwf84dTKfG5qfpLw0z0erDdAZSSzejTR64+kW
KfZ+i/wFvx9BoaU+fp9LE7tegcGfLXDWf6WP8EF/Y45OkrD3Itnx3hoFD2eGWEIKRG0GwrbJoCMK
UoXSrOKrNeKJpERLtyOTrjf6NKMoeO77vfJJXGgV9jf8ysI2mvHAwHOzNO/F/JmyVLaXeTT+0hmg
AVHSoUf65hfiCrbBvh/g26YzIQvt7hKFIclAg29l77UKzplvFHNDHoYRX1j+3ebzDDksRPJYXmYH
I7RanPg87kvffwFFlNiGOzUOQyN7yNWWugXNruUWM2ZLsNwabxR2E8rlLA1+oqEWeNLd1aZRJxNr
D6mDgxOuQXAzh3Nn5HRX7TX81FdpkU1VQCSuSHlUVggIa0ySpwlhTcUAs0vpw89utNs6vpfo/TSh
QwL0AejmF3uuMlruNfA32eQ2QRxw7QDbutmNxgP9JjhtKYJaZ0Ee0cjk3LlifX09uPmRqe7RczJT
sNnXxqlwNi3wUDov3pkz+o1m23s9BaDihiUKBaovoZ4ludGGygzL6s6V8slzhtK/l2XHGaR3qoU6
1XmNBTbgWu0JKvZU7Tcg8KEZ/Z8/+b6MlszIEKaD/eryq3LdTww7NGrC53LnUUp4Ksm4a9xBp9Wf
SO5oo4acWNgD43SKj8X+3OQ9v0htQM9/yPEfV5Aefo44x416hMIRS2deTyCa/4l8AFg7hvRw31zT
T8mpmq5Vxa4pJN20M1Eq4X9zpBU/hDLBZBmX0us2ir2EFi1k3UPwxTYfSRi1Y5+xnOvATjlBMs71
cI5RyyyJMbu7+aOtUCa0DJrHND0RTNUPbHwS5BW1lmjpU462HQzr+t1mcu/LegFU9u0tGtkS9UO3
+gjM8QVDJRFMUBbshfrDsL/VLtt9lACyUD6uvSq3qFMRZrAD2maMYvRAlp9NYSOAeRGn0JIhzjzL
R3NIwn7pmZ5I0XAN5Uaa0ohDaXXPI/S0l0HjzZCB2xjO28eyNRrUzeQDEh+OdzXKILTTi4oeR4Iw
YlnbV6NKR2z0SeapcKBlbLzcv5g728bBxkSA1awAqYmii11urY2/btLu5l6452jlqGg9qdVU4TcF
Yj3/tm80L950n+0cbaKSdHIUFjn+WbAmqfFKUDunqLix8OmazT8dORaMHp0zIzCifZLX9fYROfWC
S83M8YxWkqD60A7PlHGaSMZ4F1krjZMD5tIveD3hY9xooSlZCL9QCjS7FSBzO+TJixxn6hp/Dwvt
RVvFWaNvMM3daOuNlomMEOpg7WIYFEaHzIp+fQAE/HC6zsZM1g3hvCO3dJinkBfDeFsxXarp1tq9
bHzRPw1SYQSAPrkkv7S6iYkgk59IOh3Q/ZbqST/gzyGv0gj5qtRALzWHIqC+C6f4M+mGIiFC9/JG
l7V7sZ7jsKGp2AZ9oDfnKKeIllBmZNDVLEU3VgjMFc11q0JVKCU5dBlADpKdL+UN9ThHGSH37GcX
B68q6f0cFcLg9iI002N+yJYUvIHwakreJS2GUssriEtG/AsW1+xfnN423mK4wTgWjWnQF0s+dBVK
UOeSp/6OTv4MaTD0RnSA7S9bDP1165soYMSvT2Eakn90MegcVozSRUuEOT1vYajGfiaCobGoYcXc
xbsi7nrVkLki6MRezwVP4mCPA2XBwhEXaA0ScEUhv2Z9DmrjLNkIdVCtu+qg7YHZs47EG49vprGw
TvMcTByNAlQc4JcJPIhD9AINcU84G06j8R/z0Hm/Fpejh9CzO02zar3Zzu8/Gsv/jQwDgn/qHrVh
Hrtdjwd2lw0Ke5HyZKtG/3m0N67tEXaGyPWEpQrtA/F0vsb9ZRB+P35mkaH0aZtoqnZrCdCmpT6/
DCGc8bBRwNXzlKUvSpT2IrjYROapdSioSQ+VkGYc9JG/7lzNv4CVJ6FXCu7q3NsFPf7RXlrxCI66
egTVAMP9/GBTD/AQPyNuD7xaM4IlUoGxfEFavBX2nhV0UwJF2FVXbv23ylwnxpSi+iJN9CFnGkDm
6RXGLfbtxizsYKnggFTlWmZCcKYnVciTfTqb+YITb+Uh5l4C8szZmP8B39XLAY4QV63QNxbGn2M8
a6b+ttrJqY2c5dTKbpl51YQzhkDM0pVNn3i4tJvXb+hP80OlYOoEqhFqsAv16hJdaQSyWXWvZKey
tkS0eosYYuiwgp2cs7bVXZrTmmscJ6GaZded91Dd4TXrcvBsfNWcK3qA+0vW8UQhx3eBB4Xh47q3
Nl+gx8PbkXaS5NIomulItho4wCOWd+tfl/KPJaVRwObMwTOp/KFojikWhSNxbAbOgCCyKVNaKQma
UWvqoGOCz96dG5SlWNaen87hIUcPe3LAgqpWHoFEAsC2NjOFKbNSjRsnoyzV49f7PUPjexJS8U+T
MWIUlB353MDSmVWHWOgwhM/TUEm+Sq2IexyQ5W974Re/IiJ6HI7EDzSyFuPjoUg18EiHCj3ZM9y6
rw553iaQF5BCXm7opszzBQGDLUY8nVEKAXzht6EoCboLbkVr6/QZD9Rh4xDQzEN+o2urGk6m6rEo
pqAiveMzpE4AWrRYG1C5bysFNN3SJjIv4AhufiPaiCF+a+Q0RoHnenj/GcWzhgNyE7Wf3mRgZEs/
li02Bt08DJgSwbpZDEjigAskKnVdhdzfr+9gwD0wIpn6qF/4ya3b+NT0wYMFB84q1WVdGvLjOZ/M
/siOKPf79oNxCRY51bkGNYlN1bOIblnVRkwPV59TYcalXf2HgKv+GrnQI2gIljqgcdYaCvKnTK0Q
wnlmwIRCfR2koM95RtEPNv4FdgaHdccLMDKqmR+PMN/rJ2fZFkkeYD6WbAuyN1nBhxZD6ZQVVjw1
knOK2UnAS7e9Q1XNb3WLOl1WhP861SzMfQvAwBi9LOLInF2zba5Re7J7wqWDBSmonSM2wWWA1xmw
Nwg2VIMJZhLe93CnECiE6OT8YabfPlR+kJnu5R64y9m81Orgt5wu1cZGcw1MLKrTOkjYa83W1EKj
qgGc2yhsCeyQciVl/F2D8vg8wlNVmIfQ++o9FQWgsfB6LNnZjyVDDbAmmGvEscntplRd02Fvo2I3
rbFtL8Nk/KXe+qMs+Ktx3/WwTkEXVANJDKtbexsA1KaJMZxY/L3/Iy6M//h82TlDYwMkjwn0vLFG
VbSVC9CMe8u08UuDBrMlaZVRDdwKVM9gxss+G/1hOoDCWUnLGefEHJkQD5iP+/2EXxlqqPM+PfQO
6zzI1ibwOzAIZgGMBuRpoCXFf/L25Chz3J5ivV08EwsOkbP9ve3CC5B46fOR024KtjBOFO32PdZk
sog/Un7dCRBuTOANioG+MFvAT+TQpO6IYe4OSEMEBoH8Ov075LAHOCpLvYjR1C7qiPw7EfC2WjYb
t9MXFJWGfTK3a+DFO56Z1Y2qRPDhyebuZwq94n+cmZY8geei2CEXV4T6xeEPVuWU1DYH1CM9YUdD
NI4FEDVAaVAlCrM4wF61lUfol8qgU0w3H3FtkH9mE4A6rzwxffLKIJKT3vuchHxeeXf4lo3j5I0P
ks6tAbNSFT8HRxWwZZ7Dx++bz+wFJ3IFmdd8JNrXhSH++2sy9tX86f1eWCKELc9tUzNKmfhYMT/+
9rntP0BObpFyIJW9WBJezmpZli+IhOYDh4YGQCLNPKWcfyQdCUKwbh2NQ5nwo46rNxlbo1p5t7F4
40r0brmoOotrBRnNtGt0k8FmazeqdmLSvIi81NwIUcLi62KqaPXkqSPA4TZIyZJLYpIZzgkYP2bu
2f21p2HrdXIBrH1BsxvJBDjNVLuB6s7yHNarRcXDxXfZ/i7y28LgiFYgCPQ8yVPbJURS1pFqy1HS
57wmlsini0K7mHc3o5HVSlVc8zxZGqKAdIgpi4NWiF1RJPwB4LgSwi3r4zdq0bgwPiIEEw6TVQkZ
L/sxIScTz5z7PyQZJzp7tE6qwO4btkH065zLvlPVj37335Q5+zYGpkREB2sBaG/3Hm9C/z7pAuA1
mrQbbndFu1v74hFo7Xv2GSPREva8oGSPjeHLOHb6T+cbHWqLrytRnIHmSmbE2r8d2ac7fAfCF/nX
FO10Clb0f8yLSsH0oUEhvTijuk4dCdBjguHiLrO5k0XPsOF+rrYyZEzEe+m91FGmM92/jsNx95uV
q9l62iiUDvv2Fnj5Iajjyt6HEYF4uw7T+/5c6D/M2yoMvPaor1aeScrZEt38/jr5Quz3si/2x3rH
5wKfhBuMFEirERofuD9harkHjn4goPEYteR6aHokvGBJoACcjtbL37NJQUJusjV75zfo1I2JQfWL
D+ApvxjWBE4WTLn8Wv4LTpoVLHp8++uQw0p8D6RCX2ftQMyerxT709AoBPoGYvyb/bw8b7L5tRgY
MCQfZIXmKPGQRgR0S3NfjFtVMTeBl3l9i23BBL5trSCzmFUTJYknH+NqUAosdkgWA0+0ckmcJQ53
hV4GWpWJS1D34x1Jupbf972i1Sf2SOV1THLUJqY46Un3i96zU0PzwGq19bIANw05saF59zFX/tWE
MkgL/KF59sOT3beM3BdFfFk3FY/yaFLpgeGuDR197Ewyrdw9Tchef/tn1Q9ozvlRG0yGDFtwxtQj
pSbpnL+yWXVlJ5Yasp+aD4TUL8pgfTrz2ABxj/spmtUwyazsM22jOG3J3FayrGZsLhw7sooucLTd
M+hCPmq+Hmho0liI7SS52P5jNx9Hf5ely5JCpR7dnvo3WvBVU1Y/f5uX5LG8tbizwRaGOtD2cX5+
KzG+BCCtjYwd/id3fjrJnlrNcL2gsBBJeOrMiWthkBSGku6zAxxCbw7e7D5exJK4nbP5fGg6z2lq
7blWwOegQtIiKt7jckiryVoz050OqicQ1T7eMMC/XByjkQFudE2hXV3hEVBZwCpsJhI+6xLePouI
pWRklbqF7MzEvunZlL6IroIwaL6nZw7kCqyaKh5eDtIsCWpDLZuxJK42awZA62i34L+eKIZn4T0p
lzIenCl9ZECbfc16OSD1O2GVw1Rj+ph9so9bhCK6e1ZOukaql9iLACJ+bDG/mKyvq/2Lbo8dgVJS
4nD+Jq3gAuEeiDz1XmdmoCn5zd3gfdkZC1KiNThA4Ak+YVmZ4OAcbSLEfXxTs9jH0BOyUcT0pf4K
/VUd67vie08yGRFOthfI7n6nCw674IF7tQTJIMSu+KQfSh4IY8FQ6eYp4+m9Xg9N+Hip3Yq6NvcX
Cfae0tTPoOOdtbGrnuKZUl0t0tWySJJIdqZwI4JkLAhY40JsKg7khO+/tZgKbhmgM30rhLyxgGwg
n8cBntKRB+0P3T0K3EyEOziYKiRAvUG5apjBMgd99kI0rt6KeYyhY/t6me2WwlI9BwCyj6kjMwy7
bgqkJVyFvg7ypf2Y8YrayT24lMjLkEtrZ/FrXFc7I8c536Mn6+WUut8m/K0uFI0O2kcyZ03Roeei
MqF0XnuU04N1vskBFmcEM8ogs6FigGSvyp67rjPkjwfSRx21WAPj3N4xV/wINSQF3XROAS8VAhYb
zQJXmoQAaDK74fzZziYHVTevE9R0D+moTBP5+mEZafVxZIZXjtG0IEMY1/JBWlay9QgrP+Y+aMVS
yCYKZXTSQavLTCrhOHJwGoSn+fXLdFYTSlc8rmFOrBDl33xqr/xTAGqV41O6IwGkfbe+Z1lWlTlw
1i6lnVv9x4WFR7srPi00X27kZ3H1UHt56r/sgabqHg3OQPZwPITAtUODssJbcKnyJ+BQr2qksfVK
woyi8nLRKEQgdtgOEWLTmqi969a2I2wlYMbwmQNR6NzQ+seZjWf1RSYE+eRtd8c8MGI/zuhXRIy5
W5tAdL4vCv+lGl160PFJ2xvn9VkaBbj3X81AjAi2TR6rO2eXwjk1WW8CXjoy1b4zrWCANlzoK6vp
jAm9EGhXS2Bhf8gBd9jYrKZV4m/l66IWTdF1SGNWV8kZJcf8luf+8Ky8wAV9s/vfaOJy6PLQgmQq
RAFozCP2S9kVGHy/VFn9CuGzNMBKs02RDe2W+GX7wSFbADFXxV9w1TQJUGxFU7sYcR+aXE0NzjDp
KcwLlsMh48t2D6SiI4zseNIOVK/mDw8LB3AdQmPWCp37PYQOfJbzvVifucg/ZLhYSrQjh1MerGBQ
PE86DUmLoD+QLQcv1bwDSMyEkMZKWM8Sihle5f/hTEPdS8mPPprkb3cr7dGf5vxwWv0j8A7L7UXL
l1r+TNWYsLblCC7ghaFenOXT8lNp2TLfEC9niO9oUKUpC4rOzsYBsNZe5S2cUk53ojVK2IMzEZnU
sVTZfGteEJOkntsCI9nFsgSsGw4Nf23G463RtIkdfsEp1K5PoxHzCxCZz5ffbV1DW93qVFvXncvL
dIcqJ9S1az3asOvb5EtAnaXgbTy4Z3NQYsHUgqaHmU+BYYpntlEW61D9Pp7cQ6d0SoRpJ6f5NScE
TlB55lgjt3W27oKR/DyD9CNsFlRKuqfOaaZHOzBH9J64OVPOBW6EXGwHAv2+PXxQD7lftttSpzXH
5mGPoQiBvkQZGWPanE/Up3pmT6pATaVczUsfGq8PGYUOOjtmkMzKSTwxKaXzOBITxsovpuXxORxE
KWYNUL4o9jx2ZmnlIxzr3cHaQWVsT7WQskClHuLp55dAbjYlipzRhOKYVmaJ2AkYCVTly1C/0qqr
7q66KRo1ebMgVbh+HB856Ht8CiPmGgRL+t8NVJgW5smrLsNHYgvR9C4l0MgV6rvO2RQUahAlPqGf
9hnCTAy+7abxaTGmrsIBQaR/XodQXMXmTKSh8WesDolaL1VvYGUU7xxzPKLiBUByYnnEfPd0Vr2G
1HoGVDBAFT4Ub8lwIVf2tWzSHP/+pHECpcFHgr8eWj7bwHB5dvgIxQOFs9+N/qHB8r2ZOxNOqJ76
UFDKbCL8zYHLUEqtbjrIezB9KlEDrqsYe0vaMhhhSDVnbOskMYCen36k0/XhkLA7kx5KGFPMynHY
DNOHYmeGL83TeaGpy8EoOchhqhPRjC7AzDCopRNh3ppHhU1NDBK0SrBlFgkDSgCT0LYHkFBu6SFX
Nwyp1I9WNarSFMuSYKNqDqNMxR0+d7q0CCPEreDXmdmiQNgyAe9JUs2Ndm7sqKQaiFdZvoFWInbA
TTr5Rs7UAFUlu9UQyVmiDpb91iHFhj+MhQOoWMaXK00QVT89WRrpSdZfepkvxdUc8oJ1B14B5X2L
A12t88JSBszcHI6u77XP9TDWxOHRj+Z2CMZ/Eg1mUDiA/wCTaVaK/Le7zFB4/R7BDbVteFFp+BNr
rSoU0wLFKmgHnn2xP7+GZjYNzige2HwJ3WpPW80w7Jwna5Ve73OcTUBYvAvI/MPSE9etIq3Eq3qb
wj3qt1+PlEGC3gVFZ/vJTGDFElVhqBSMH9v9rAl5sUaC8hOqdBd9kMVsSUJWjmkJN+ZpkdL3ZMJk
tKhpYWkYWNZdTx9i9IvezRwePk7w/jR3UBUrE2PiBerADFsMr9MlzCPtxzPhKhMbgcq4pp7KpNEj
DEkEUZqupXDKGoO85fgLGmHzkrGbugDmeYobhSDX3++7lhw+EtPQhaBFW+uYU84831YLzjp+qCXu
qqtEaRAePRte9pZc7Va1qi+ePSgs+SJeBnmAAtW3DtpPwuULY07UK1CGJkBVGtFQMNxXkGtekPt9
jEgsqJ44m2G8d+NvW/ZECHzzsDQUlNAkHdExEI0oecvxhl7IY40q7yb9EzjIv0uuLtVRRYIitlPI
k8oGzgaaOWltKuZ/JXflG5YCr1CPM4YkD47fFj0xG/MlhtPuUBP5daLqGLBd56NYXxRkgZVFOWO1
XFfpQqmaJdBmptH0vM1aouBtJ0rGSZ11v0IPA5VmyEN5dPjPlJJOJkle5+zJ7Ghtk9jliLg11Ft6
uLV508I4IDbHYgq5WbpcXcmtCjUbGk3b3f47JLR0635Q9/MPeebvgXt7A/G+9GOGbMQKFeaRKGT8
JbdQm7so09k7SLehoijuLu6gzz+M473SO0Dd6Hr0XfY15uDYN2cipTq1CICQi7eMxN0pF4ufma7z
tSdnRtyAPimAaGxlI4NJsqTxk2eXJ02RutqkNHGanybtaLuBFsYmIUva2VOATwUB/m8PPT/RKbTa
nR/NYLpHLeJscVuOpBNduUwt0uzrUkxjKdlG/BygohWnQI10CGNGg+s5A7t3m5DDXpfc4byLK7U2
1spP8SDFFmIvSwcuqM2ismFHfvkp5Tk6uLYf8uAaFKNGVwZeOtZc5by962iWkoqI2pdDnatAPQ08
sa9Gr+XEzUQn7LfqkjdximrLiLuKdugMRtLOca5InW6FsxmQi9mpYjzIVztIG3MKZGF4s1LFUBId
Z+mnsEWN7NEMUV7dPO4LYu5Ih9U7nyOJ117TJGo17HLPS4Tv+yqjXK5X3uQ5iWvrc9bc3rCiQXp8
IrkY8xvWflHCL6/PnWWS0MR4ZAqq+gyQCHyuYY8FMwx3PxCwzX8nXnDBYvzSSew45Eixb8edjKHq
twj9UqyzR2zirpgMaWnIvWjFrK05zXErvHO8J69o5J+XAM+aAdbsm6VuvRljNRnLK3dkrfuFVTUr
NUR4tuy0HR1D82WGgF0llBRTOx4mz4mpMhqMXEwGppjee0x11Gp4Ot62Ya30PFDygePJiTwzJ1Wv
7bUxDNudTU2e8W+hA6H4eQ2GKpWs47h5ac3dKvyx9vUquecmCKxQPYJ6fKMx1Cp6S/R4AWc56QwP
+d356xHTu8b9BhQ4RlXucw5jt3WwgmZX2JqGrF6L6BkTlfh8DJqIjY+NEw0h59qtR7sNEi0CE9Fe
BjxGcIQIL9YW6k+K+1cf/KML6cC45GjALbbGwjPceHEFvfNcO9L0ieVgKFOyjZvEabwiA6c91jVP
pmHd2gdWyMQ5X0cOjmpO5UF1ZvK18Jy1gYLAKr6q50qLjynpp160hcxpEUWqT7het/vWqs6OchkM
UsxGMfRkwEZoOSkXiKkfPJVpxl4HBlBIwLUkbSHi0hVy05B0P3uYCvMPrTGJCvM4oAzKQ7lXdwcQ
nN4jPk9MsJguQWOtgfxdyreDKlRN9GdY615s7jP+zaYO2c1z+KAwflV12Egww/QHjig/ydXwdNsi
/qnUdclv1ySOB7fM5TABqQYVRm0qCK9OjqX4TkiStRiliLR5bB+B5YPfWkT5FBDOw1rbUAHXRgk4
x2yBVme/aXkGR7KL4FfB1lwVH8W2vZ2Y7sJcgzyVTNfyLKW7KDAlamOmdw9S868Y02RJ0Ko+A3l4
uWAko/OG/tGIKegNnedk7KmHpcTtTbGt1PZEmR2FALOMo6CkvdjOOHDw54DyV+TmwqV5UdS/Z4IE
BdnEJUVhgqIGxq3Ih2B44E6F9N+lwfn8z0uu/5EvJSp7k5mStlJiySAr5eXzM89YScfYJ9py1aD3
9Jlk/PZ6bF098uiIyTbvqgz2avLhopuvJq8P0Gz37aum5KYmrn6d1fYmfGAT/ZuYN4qj6YZjV+4h
sKNAPANIcKC4FqnWdAgeq5NQw+/IIZb2AoEq/iFRH+RlycmKCu1567yDXXwsLo/xF+zvbTucr0gn
aAgBOAvv03PaCC8H4Z8dIOdUxIAxKkhwmOoonGyuv9HqqSvb/QWO0gaCMb7BIT+x4EiJFs7ZV5+f
LVoaECh+UW/RIdNEhyeTmV2L1WiX+5M/B5DHvR+hru1VRA0CyS5xHLYutpaTft6dhXHnpFjaxAR6
ygMnzD/TErWQa8mOGQn+Ie8x7mhhe0r1MywQv8WIqvdty5ZxwK45l1HCAvy01zDlsaAWCR6k1u5n
BFGBs/6xAMCovI0A6M+scnRiQf84sYab6Mps89nljtPzX56zNusnVkT6qqUnQphgJ2ARo9po4O+C
YEXTaj96KMWvJON9vzJ2i7BIOvR9jCsn31TUcDcmnFnj+3HottOoAGKufB63baDBILqMGXrQcYo7
sGEneDLnC2DIFxzki3q9sbVr41CNzcapOLdMjdYyNm6q2E3ssoOEVXbmoqArvD5J1E0tGydaiHLK
BkhNqTcudtCQ0WAJNacH0J+CfBNkcC9u5RdLlOXw/484I0GydchYplXfN03Kt2regPYWec6KVK54
RD3Y1v13VCYk9Qs4jDU7WnK66NdOfKM33iQBOUCu8PdOXOFCiyFBSQtHvXAxt/xJjiqE1aVqIeHW
IZxgZwl0ptHN4kg3Rx72RA2wCtNA8jHoSt2+c2+34hzkuSLa4pf6j3RFk7bLgO6yaJJgc7xd4Dfv
ONVhL/As5DMVm1SQIFLJ6lUs2VhOvA5fy4k3p+c6DLBL2c6PGcZ7PN1tocaxYNLQeKFE3/rvKseU
JcLVTJShLEIjZLy8EQ4OVItjNiNE7sE+KYPqWW4vH0XDVIuUPpLhW18yeI+l9Gwn2mRmKbANlI8z
7d6q+GRt+/Wc3rFc514F3sjfgu3TUBDjQqAOohOBVAqI4AT6JFvuAFvtXnRCZw3nIk77xoSt4csu
b6VUPMIoYnkElXXoPKSzZ8/8sToWpfyZJFixgYqHHsNrRHg29Vv01iLhetPSHWSvYW3eoOd6gw53
CpAHppyVabAqcWSaVFmJyrdZqQAeakgcbFH3JlmzMgwIC3LEHjb1hc2Cwf/voJsst/ec4veVcVSR
bCU1xEo06FvTrDq9ePBTLb/Qd/2hFGJOaDUZyP34Z27cQGKYfXStaCU7ZE2E/tfKBaEOdZj9XF5I
x2mpBvV8Yu9TKOzljpfNbnf8t1jkJFZ1xx9RG/ibvEK59VNkZO96bGwpGM2cNj5chPAWmjF2Y8uY
rSRKVUNn5Ui0dK2hUN0Ogagc3e949Rl3djGKjH1YojUYV9yKsKxhqZGDWAdqnQQKIgUwlnxBYugf
5KYh9me0hOrKyWfCbLH6TC2InecVtgZRMYbaVq/2chxfSAKDOcfSPyrVVA+nHd5groRWoZt6gRzG
JzalFyXD7QPTfsELMkYbBL2PORPcJXieKZR2jr68+erVO7bZXKePIURWxvJc/vTVcM2993UWy6Gq
hmMR8AtC/hXmyt5iZFzMjFjRa+sr7IGC9k967twXFV7bWXZKNKSJnnpL8xc0o5Mg0M9BCZWHsYv6
tLGmevQIoDEg3ozJaWOzySu21Q8pcH4O7wmMpWQRchC2Sazxd0wOFg+381107/vakZ0gvGKBzE8s
9P4EVKwAAvnWp6Mj+FkD1DKSKYrbhOEe00suMraILNo/9u9dVdTT2AI/TG61jEaCIAvXFLRFToUi
4Y9Ko5Bvxo2l/TFuH/uVArXya9Js/k8GbzoYE+plfArvzVU0sghzMh+aYSz9tB6KAWCKrAA+ZOPo
pfWHubTvsL+qchqDqSAg4WG60N9MOTFJbLyHa0B7trctXfNWUvNoFNvo7u0EoLuaRyI5noNPriZy
RkTngbkQkPwABRS2ZaGa2PH1fygYAjI7kddANIZ6q7i5yjcaxPpFpUhlk9z5cSlleQ0/El9odlZ3
xeQpjtI6yvF3ARJ0NhA4KhefXqGPUSGdPZiPADnh5uBYJcL6TktKf+k+vQKTlSExV58de4MGQNXF
0j0pbbJTG/PUT3P8zI0uS7tfH+67XzwUdbrHkYuvRx0lfpnRh52xzK050mR2WNLcc28WhaYpUriO
dvfgYbtxV28Lb2cBg+LQwBzqPlbV3SDR4z7gGWASpfSnn8XNtha1PESRINAElHEqZMOJryZqL6Gs
EJq0vgdnNo/hHCNgBBb4yX2Thj4JQQjw9PipKHtCzGzIf1levOVjvKQ6He96S0iW35rhxSX6Zr13
gOyXTwYxLbMsgWYCgjDeanh6od4YQtOVkhggEUV8qXs0soRcAcqvpGaFvyIbLWf0ujlGiadGOhX+
I9cY73K2x2k6TIbJdfsX9AXb1HUyIAdHLlnEeFt+bS4zMnaN9rjagyEwrCYC6eENr7/fQaE6hf1r
AwAjqDGD3GDASCtAjfkjXbnmuxd5un0H94J7k5oSpwxO/KIE68/AAJY/e7XHVOZYzQyVfHWJCgj+
h6AZZ/UuFRmc8yU2SYreyQK/IWndK3gpeVEsKSFi2w9Al2NGTwQsIQpMuosSItzk0/Ziewjvd0tU
QFjeDeyXrW0hrHNjU6Rbvt3RllSWyOAeKNesGuuU7SpGGvWByDk7hxFYRIbOfUfLMlIhgZtNkxc2
vmeYV/LeJc8dMI9Ei8ZQPnYkMZU3oJv6bxBiUQ+u4ujM3CSjPohZVJWbjC+LF3SBSnTRrS5SNj3/
+64AH7PU1msEYcEkJQE331pzBEl1AlYe8fxEc1CbK+5KfnJ22Q3CNho18/U2b/juPzg8kiZJv0Ga
Qd4LwVQDDpHEtyceIXQZwfKOR4otc7fIHO5YHlpwLxgzAOAFDiPgp92mqnHbeL9r5h5JwvmInP4X
ZT3EDpPVPd7R0Y5SuPl3UtB8dJW2UrF2KgOHrnrXPhhkDNmtEsI+WzKZG9uLf1U2fLHP/fXPnEVv
Du8B1YsET9XGJBWEwo//qp3qNXRgaFD/mKR+OolE88FtwThOzt8OGdcC2hBDWBtskOgjwG3aT1jg
R0d5/3LG/53p60yOnjgx7a9gs5H09tV17L3EXannBnJETAL4oVyTjbDi1uRJCiEdfc4uAb922XpQ
ADtiopDlA3iXh36uK+SXhLvdJmUgwtdxylMz97eXLA2RIyK1uokKiTkSkhK8MhPOZBHcfKycuXxT
TV21BhcdjUhq0MEmzrhXyoOpIrmiB0w0aCoYqa+qXEQWDbDOyy4DqG4Pms9wf41SV+nFIcQMC+Fs
2KL6RF8rYPViIp4bWOXUzEEjRGM9JQIYd+ePSWjlmO1I/d8shyTn1NWjebO/D7/pLUyPe349raAH
/LUA9sLLO1ZZ55GN7s6Ot8RzhQ0g3ams9sIMxTPqaNJRA9Ny5K4gxHKDh3N+lxXKW2aKEl4t40Xn
xnVo3ER7nh80C+01HE60me0e0HJcEXGzS33gcz1qn0ugz4iIhWxGROKvpQMUYbOCxHrqTmoVaxP0
FGZ2D4kDKJZ4+l9xPnwIATAD6e0larqFVe3gX1XlsIirgxa+sdSUy4k2jKMOvdd9GliTPEmiONiM
uuBIb8EWEfFaAxUAhRBLPnShPNDQuHpqFn9K/yowl+Nl5uqV0NPkWR1/OUPDaR+kRnbkCFScJCNR
iNOgCC/TwsYQN1tYoLLstPzyww6JI5meuE41BLujx8m2TsmlC2ZoR8LjF1IctBHeoz1u9HUpkMM+
ZyaUORvs8FKJFjBrGcWJO++rXCEr4q5PEZh74Wj64KVjXdEY8V0op1ETuJs+//IDpQs133m1uXy5
N3c16S5DxEW+iixxeEnR2Nwgyigw43ShcM23Hcytk2apfPOWLV9dxd3GW+MqwbPJCoKj+6RfbzG+
eqrcrVllq+W1nDO7TgcjEFTpkgBgVM/xLmXKfpUf7rBUszHjooBfmYASuGul0m7COZGZ2T//IvZW
n2VNoFR84WsSHeB6zhruFtZsya3Bws614XbWRd82KPD/u9i4k+o38mXZ/TPJ+Msspr78B0wZAKfb
9Mb9s+z+GacvmZtGbci5btfwIuK3oTBisiZlMNTbLHMeyev6f81+gpzl+ht0V3UGMeRl94vqCEf/
KZzOPpR44cVJa/vG6rgIu0Hxv3QVwaMut2tvDef+6j/UdsosWl5XCtUe3B/xdrMSr640siq73SCX
jkAcO2idWTfOvbHqR2AhlkK/BrkKpDK6TscDJA8WWqTbbl3eOtjOUFkdSjxvPaR1LGiad1O+vWjO
/DU9IprN1d8DzQ43t7qzovmURgbQpV98DDKVFIrUrSjLJj+mM1Y6sJcWNuPid9FN5MVVZg7cE1QP
vRnCvFntFxV+bB+baVbfhZIX/pEfiyckG2faJr6rE90D5n/VA+P5cV5TB+CPkPpCHeiysjmGAVBB
lu2gZpIIpZx0U3yRcdv+EsfAjkYi5d7qVGkDjCIqBUwWAbhsORRaWifshFeMzUNyPV6/scZSpWQY
ii9M6GqoXaUs59uCt3OCMFP/W43qUIA5NJHnubBbb3a9DG1sHzOoUDzlv3AmIxntXsgyXx2nKUAa
AXt1CZrG6OXACfL/7+KHJ4/RLMKfI/XvS7BE0hZ710+mhwl7Okhe+uQnSfclk5ZTo7A27671Ctcd
8BSwtNGtpP+q6k7aA4esH3MHEcVc0TA3mxb/+cwRX92gr7BOVbwzyfG8rdqppWOnX8BBYmOJ6gB1
PhHDOkKU1raaGRs/65xxEhQNYfzYRp/XfeX01qMDzSxp9DF5UCE29HK3DyVSJZ+f0uciBqtzRtrk
xBxah2asCFzxnmz5b0CKbx4CfP6Kg3CNrKhyEWAK+0LxIxQyh6F5yLGC//Y/cUFX28tUJiQn6mZr
MEY7r/wYflfGwBCyZc1tQm/jMRmJG6aTB5vkKevPCtN1gEjLR2Z0w8oZGE1sYJAP8s6u9F113l58
nLfMnWtsRkLnMIoQcd7DukVFpZ3ZgQKcnJtdkgUEJ7TorRmVuQJgaklMFfgLU8nWH78/EcNq6S+Y
7yzIGJ7JGhZ4yR1+9oMBAAO8hIqSedFXwY1xUU9wXTUuYD9j0jvhjlEdl2mV11dp89Prdb46AlCM
Xwj46KZHKw6KE7mtTY3FDEEeWFJiMzZDa/HrQrMCDl52o7HCGYDZxmTGqEgYff1P136rBDX3PTSN
/tdDhSLQlyCkUcUKA/WVCcnP/9jLDtnKZYdH9D3Uh42tE9O+6pCxxZTjrUUQi91BGaugFsXFicDx
Xpz2Gk6fRBHQEFNrexqDHdpLYPcvE5HDmaKH6elP+JLtNVhLFRMIT3MromqiVAHl8tmRVz/lzkWW
d9Uvda9C11tTRAgreS2tYtosVuudgx/+K39FV3WeInlhvqHAKXWRAm3VoIQRk9wwBKqyKSpqz2IN
JLEjgqEaenC71Df3/Qy3hpb2+iZ6EElIYDKmAfnE8LM4+MqNj6Rt9pTQr67VlcyiU+35UY6mGlq7
GETI0VkfKpGdiduVYizlgAakAQV549HyVfCbqEJUt5BmsbcibotTid9/NurtSVsv2mW3PVuYPd7i
NaV5zfslrWt1g+teCZO4SKyzojMSpCUsV29ThwxIv+7nBFQfjXmvfhqJa4rbkpQZSewXO7WFhEP+
bK5uZUiHP2/fNNy35L11/7j3Gx6XVpa2jq4jTNnikxTe9ixo6bDNYEyt3RbDKiU/O1B3Nr6l3fLb
U47iBBLpSTMlEYFbKtXt6BEefSjVktv8wizhPvjXExsl5kOrRO72QoLpy+VxpXUfLih8urnEiELo
FRttk4aA3Il5zvre5AwMMbKH1Zpv152C1BdunI0fKkpWy+OditPODLd3RtFNUewKApW5o1yMQGxg
z54cGG6J961VpMwl2VAzCRRVq1HUs1KxuMZbtbqjBUyQdatp89xFVG60ysGIXKVa3RrTESlZTbCU
Dgdu3Ftz91+ulvV9VmVJOdqs/2zS754Hr3l/uPpA265QDhfusVFU8mLVeJx9+rooJNqtquaaykSd
5UeA66NUpwXm06VnyMUIeiDjdVtnxgV9eLvFzNzDPSp87o2SXoh3yONnRIIs1IO0gdlslQ+nN08i
/hmJZtDm1TOm5MCs+kD43zcY2iiBj5Mfru0ZgX98fMES5+1PEJKnRZNdG1qpsrKGlGVOUQVserhg
A541+C81yIHIOI0FELlabWCHsOBZxAW8l251VJYF+JlW/OjwJpDaRpo3vU1XaokP2vxbN5x9w2t8
2taxYYEBoCogYlluCbsmwuFBGD3yrgmzBzXrb0CDsKo/QvZB4Ta9rUUerMe6xqJb6OYl8N7KtWX3
Os9ShRKaKNeImGrmH+z7n1SdIf7rmSswSuV7bDfewV+XG7YW1iGlEKeXk6Y+Cquz0I9QDxOnKk2X
+Z+PPGu/ksTHk9VJqyVdoQQxaTBM7XJgIjfA/rROtj8ImMqJrREb1s/b35Cq69nzNtB8g/yA2PuK
NqFKxz9KhUTlKa1odvYvVefLeWEXp4YBr0x280VkcXp4LQwUH2uoJflMOk48+IGEMZPZck7Ywb92
KmubHEC8UFvfaX8dlqQ2XZnAHYKSbM/LBgMr4WRmdtVhinqdiDVRynOKE3wsZSKKMUEZduX10mPg
4SbSx46abVea7iN3bXDNEmLNlPPkuI6Q7+U2ROhhpJ4RbNdMLXU2JJdbjZ6GokC2b189FEtmq+T1
14RvDEQvmAo8Q6Y1zlJdRojeIK1xmxGIKO7G5ItKGzwjfNrC64zN7NpuEtqe6fcxmA2AEB9njlp5
T2QgsL0heUpA2lO1/M9ke+UpiG/hLyM7P6O+iIH62ps0qyBigrXhjpsAvhTW//IqyZSNrhtIrM8L
jdym7YM07Gq6MalL44A+NrIWUKBkOXJq3sWV1p0bR3A0HAZfooii7oktKw4UUR5wLIYtR9QVhAWL
p5vjAfYATOnWPvCW/+RCwdMB6ma71HnkqTs9IqQTExz8TnqfIdwPmEQxfin1Y10glqnXP7srSLFf
AIXKiZs26Ysii9Pxmizbtx8gy6NK29OaG9eGBHZDQJeUovlTcYF6bOv1kZf+FTMiWBpHEnrY47K+
8A33VVlDkU3QsflQxZxvbO8YLBiJe48IV9h2RxJClATIzFgVaOz2aryFzSRJfxuVWhRFRWnteLqx
3vVnEdzZciQKST3idVGOMQj0jP4+g3D9b3wai34EVgRX7SUuEFt49tHshSGNXR2FIt816N1GeCaa
jg+ls/ZttSH5fsSiKGx90wq7e/cF++qVJtJFa8xi7Jn2UZcxU+oZZqSgLSNsmBjG02rWNJCmQNLs
f5ncynScvafB0DDzxSFSZ9cjnB2lkjLoRnOLELZ/CoAmhT6TxPHO/bN24ubZsB0OuMYErI7+chyO
mwCgNE+BBbVSwtpwA+Hjxvg5dashvdUnybHBfGadS+iNGsX+HxJmV64Wv6xBLsQvmcwSmv/vfQn4
FgMf/KKo7+cdsHKdmnq0bo7YuqLa8Hb2sNsUl0iDRh5E6a1y/I7FR0qzPT93etLgu9guRvn7Ka51
GdafZkjiHCQKJOsQtC01DdymPhKvcz0ibwJVFDbB01eIqqGJlH5nmfIGKiDyHbZIbR2nWnqVix6D
4pA/abiWiRAf6IBhb7LhX7dCdiVFUWOVpJMPJZXV/qDirgxHxKTBAaBmZcJguqIyxTfn8ojADf8o
r/dN/nSaO3zMWsnrNH57FeWysGdDNfSzVcw/cFC4VdLfjpF/i6CcHz6RY2Dyhv6vZFn2mKaOFsKW
LtttOeSBpG4DSq9TR3d5RwLf21KHze5MsmHZq8IeQv/JRcp2ZYC4OCNSdPOqt1KWpDivn67Ud7dQ
Sr7nC2ge2/VbUe3UnTUI1lOkJNx1q1Fi0kxngZ8OvTVbdJ1x1G6/Bm+QnfsqgRKKOetlZXg2injS
M0FWYI8z86mHRcSAmZayRtGvV+devBIW3RmMliRzWcFcBQUGz0+imEhXfMHE5mFjF/sV6AUkGZ70
mxPpoIAIO5FPu/p+KHD0do3S1sZCsZ4Et4W/wwxtv10/BWyoX3dlwetWd45S9K2u/RvTuyXcAu0Q
/cuxA+JTYJjqwpyHrHs03qfT7sBeky+HaRCo/58V39nqQUK7xZhJfTpSoZ7jX3pGhriT4RvfQfHJ
LH4cJxoi8vaYqr/7cpN/k4VeBjU7Q4CKfMAnwjK8yi4/Zod5Q/U09/SNg5rfU8F1e55+tL76THOM
R6+vJ1mzuXfVevrRcZAwzLU4KQLy/7WpGu9MV7CrGQTfsuJnUAVa0GMpg/QCaKDzq8Gbov+In1dK
Hm+WZoUfKhPv2Hc/YI7U73Bq2KYM0sZS2P4ZROXf1R8nOd7dWnSCEn3zvh3DWlb+Fdu4aLhwzis4
Y67uypS2toUhfmxnzTAfOoe0MFCcEjEPIlXBxcLc62WWj5oNZQHbt6V0JFUrLYsLNrdsX/rhN2Fw
Zic5gden67dF3P4jJJgcM9dqyLjS97NmcrPOitXrRa2XG0L89TgO4Kdm6kTC1lrSu4C3IFeAD5Kk
0qFm5HuqFTf1QUJq0nsXJMPB15VtdmkHCjoHRRGFKH+6acH8tH6S5GF2ncnATMQoI7do2qR4+dLW
CgAnKdYz7wnAhlZ243AeNRmUEPXmVknK76qK9lQIkjuwIIbKE15Fg8hRt6NiMIY9eHj0+20rnhiX
qs+RFLz0DFujTkdcxFkB4mSbIhsEH9xTqXuPdYVs7KS8fj+5sDqjPT/9v0V7kS6jISJk4QFYRgeJ
+sRxp1RyiGdsNow10HcY0CFicgtn79rXJf6irg10avZvUF9QFpU7gAMHdZiIuUUZgvEGncnuTuN8
9D474eWHZpIlkA7gc6dhv3EBjyfkDB+M/xEIKBwaSiH/DMrSLOWv6kGUQTgwhvSTwsX0IZZrKYWG
LLziClRJRDbKROd5LRUXny1ENyXP/Y6yzr9g8Gow6kGRAVHYa6lu0j7HtNQX392lbXULfU3cgGET
vnJkbnb7NTtWR5MRehEaZVBMUWJv8GMBfQlfp8X75EzR8RM5+l6I3nUNwvUZMKEr3rSfRMvCpOgM
uGUt7DCTKlElrNXioPerkhTOnMP6moRCddaI+0D8LigSxQyqPZayrgIqkYmoVOp0m7AEuUvZ9eB5
kBMxIGUapnfvSCaWzDMuWU6rsc/E9GZytH9xbJ+0Y0lC9Ka9pPqi0kfnKWJE0CAJkPvu4xlA1Xx1
rzqzjBu/jUg17Hhd5TWu6/WvkkJtQJdm1upip3ryG4e4qLgC6DaCtiwz6VReS6m6k08ovJoMUS1D
wFyQqUPRXKJdWhNlxxAed1HysPbqnDVVrCYwWW4UWs4Mv+cmX8RbCSI0QTi+qD+Wq2J1cyj837Z9
O5nKE2cctpVw/Yt/jxO82z1nGc18oqVEKvwyQH77RponBHZzUt4MgWULR2GESFamBvmfo7BCiYYK
tM0Go15+0SkvYw+paO+JguV6F/fQqeglgc8IgfA8gU0UWMvnG1PoXmz5sQ+oa4WJY8l8KNMpMc5L
8G3BuhApwJfEPnRxTKQX6soErg5+wJAIMGjsIcD9g6OrvvZ7fZQbht88xPD21R+yoD16OX43xfi0
iHOKQ6idDkRv0a7AnvlcASim+SZKFW5jvv2ZlNSUObAHMdilwsBqyNuLHqDji3xxUCw5QQL7jgRM
DQnvqpMp70+kJ0qAsj83bguYCF75svo1rQZCEtgt8DBgA2+uuJoqXTEKiIMat7D0lPdpwtoGDO3y
EPufNUTqMQSODnNK1E+Goz9Pa/YCRbPwB5rfigcREAm+z8OM9Mc5k5sCSkryko5BZEgCdyjCQ2C8
irPQupqDYhJEgT6UNRafbqQ9OVBhyrzNGBz8rmsXogiERg4dJtqzxiI63wmilDEpUkRUgen8riRT
y9Kuh85aTbOMAeS6W2BXotkrpgsBCLQPraINnrfZ0asqJW8nf48DzOzG4elz+ZK6HMt0bRGCzAqJ
oAPD3qr0DUFxq3yYS7Ogk4EYYKf6p9ZFVFj+6HGAs+m4H4MGWDBeMUVGYRx3PTihv0Px+F8n5vxO
eefcF29j+PZ9mSEphzsKqNsZsY+QgAo+Z1hYNZmUlCMdt8edUsv/KzEc5zqs6pr0i3piyIiOnuah
beqVJ5iUHjG2D1LbBAQzv4Q6Knd8+M41dgSKyKXhc1al07eTyWAzowmBJD6KNzAHLfsb9Tr++/jU
jajWD2ASBwMB54s8NeZ2nmEJ0/6qmNY4Hbo8ebjogXrwa8BtoA06tiSys4KukyPrFVFT7Fbr+pA+
+hYuA+wfOoh92542sjYs04NUpyQEFXSBGZXI9L7O4Nu1Z4/xiVVZq5VO8eVXCZd4VX9CqbkYDr78
NeA4G4QSFVhCI9Es96G1nMeqKDMCh1zgCp43c+fL2DOfk/EkghdXmrvssTzepk/RlxLf6tcK0CBW
sd7Kdybl4eOOzF6EUUMjd+G0jpTr+GToPi2u/2jHiZ9Cr7NHwax6QfdqPHYOJNNaPcWPS83o+CcZ
tW/g/Si7F9Yne/BMJdgp4M9cTNBwl4DOIDnCzCyoOz0q9CJus38D79MTBDoERtm7YSZKRZ4M9Ets
RcNrCdWOt6XpYCJWZ/Wqh2KfB88oy+K34ogxFX2K5qKxQ3korXFrJS9IQlzuHo4UtqiSqp5rq1+P
z2PJVMh10n2GrmmF2E3+GUGLXuPueenj0NUWf+9B6WvS/fKe/NMOl0GgNM9psrbAY6WkbAWkTesm
oBdUa37gRSBJmeAXVj9Sg3yx1LEpjzfydhMwgUSogDRWA9bbtPv4VA3u7+aksWyCINIZpy2d81RJ
ozBtSm0L/74klSQ/QjEFBCBK1xe4u3rxqWGwWf8sRD8xgqkrY9uZxKSVNpdRj/gARjy3ncgJ5DOG
vGY2PqqLCBZnpbg5SHuCoQmD4CwExzLLXMIVPbW31Io8IQPysPODJPxG74Idsf2C0NqiJw5Lm5X/
Gd0m87/WJANBV6pgR1GzqKtAE00W6et4QLPa9SfVfMZOmcWrS0/4lbY/bZgGJuM6n7EexNkX9NbO
Ae7x6exeCxI3OtlGIxwmTdrJ95KcUfPsnIXoKnQi0CkRmpvNIE5Eo6rBVA178Gv5+JXG65h+9Cwa
KnDyt9MRcMM9JK0ZNMQ2Wndi0V8iYMwjK4uYHR2a+YdbL9ZPRxQRuXNc0RtixTPTGw1qpDUjwSpe
04mFqhJjZUGWhFTUNt6idErsBm4UkVorrpb9HFA8mOpM0Hm2rJXIqYphKQcyndXtfwS5/EgKHWjE
ODzCVeQ9DAKidqZ5uZQMegxNpM1DwGzVxi3SvLu0senmwGlIJEzh5FOe4SEhlcnPen1eFIh8tkE4
xVW6Fwk5JiywLph9JOBcMj2GhQd1gtTkdK/QH1iWqmLKPQQkEjQUwtk5LcbJcIxW3jlRIsWCS9N8
gDxJsJiS2UDyuk6UAoi7Ic1LdshWidpOR/Jd5gulXAsxE35CVaxfAV1+1iTomn+wv2daCAfVLiJk
tI7PmpT6kPTU87LdC7+3xGds2AOkXuk7SwcNM0fXnHwvMf7QQlzLHkcDvJ89sxGuGtcTbcs5qgjR
VALesszeQW5jkJTROKTFO44iq29uMOFxDNHqzEkK15O5vGnFjTAE7uQQ1EmdLcZAzpXDq6gv3DUi
KrNHahHbnhCZrOBvk0kH6xGfPMuivNH2asbRuCSHgVVYtt/N3XUdGNqtxeGh9rVmSksH4lVFSB4R
VOeV3jcR/pz+MpUMLEZdPgrhqx0Phvny7T/P383+7/6Fm9kGrre/7Bh56VQ2W6gf/RZmVqeNco9l
Ge4cySsvNQxZUWR5igtUeUuNLImUi823/cCRAXcej/VSL4FUOxfBDsnq+HDOdgGlQfGSoTq8RbwT
inJbqyP/0MNgpN+59ERMkPKk9lZpx0cuG20TXOUVbD1g9qOifl7rX6vB9Fz1iC2zS1OafDHxTbWo
edDi7jhgIjpf/u+OHa1KEU1l2TF0z/Wbn6D4QQHMZEZV+8pI5+M/XYdI7ibJRf9Kt8VGn4G/C/Mt
Z7CSua3zseOBzvdtr7sj9Ud3HdvUS++kBvAysW2G3Gl9lTRjmA+pCp6R3BUawUn0pOnCVL3Tjfol
5v3SEnH6CoI4Bn3X7GNJcMRb1w4T+4jGMdCdiaBM8i42a2sdIGIMhfK/P0X3YAMWbXi0s0UPkvvb
EcPrsjH9sxgAE7/4BHbCllQl/E3FjV/oXhn5DMtfgSdPg699frpHVSob7oHTFWNl8+xlK1P7pxb4
1JlAVC6NH+huXBSlYnjRMB+xLv3vb7KCbxFnbgm03g50qud+0KbZL5UlKIcbpQsId2/u7bjp+fXl
e/1xaw62G/7IGQtd2kJbZF/EB9aSJL8aXDmDYlLjTHmIbqtaAw1gOB+czPq9EUV8C6Vk/DwkupwZ
6E1IbfklYimsfMgHRTy/U5sqQCGicZbtUudVNs8Hi+rsFVSv9bf1GyPYcvPAM2WVna8lThgUUkxP
Cn84L8fw1NNPxkNBGaUs3ltQUsaUM+hNRHalMQyJiEFyy4ePFGLBpHO1kS072vIzoF6OMtxBlMFV
LkfSeHrDssemUoFetUMX3RqDDp65S8GYYOVljSsK+zfbFkNZcWoXUf07N5pVRxld/uO0DlwYmFt+
rTmgtMvWYUMKupvGdShrqeoYhVGLhyQV7y6iN3uLU/AlJ2jDmvw7G3YQoQVzOjHyz74aRBckdA0r
vLypNErwww8wezsf9D9y8J2fy3+2OYl9vEWJVM840Z7Htj/jkM5cPzDrYCLjk3ntXTndxsQpYTuA
QRBVUMMo5CFGRuCDQX1j+LjIj8APuu0sEUyZfDRdDLd2RbAQAknrnd4RsQSodLupxbB/J6hJaGu9
XQO3uepW49gdFjCey2DO3CExhQIAcebjQN6YKWTLOrpVDTGd+jU5RzBvq8CU+ZGna8pWLvRPbhLp
aglDEtPar+apUQypkwrdCtyAKy8VF1yu9kp1yCHMrPmb0QJUxiEmHEfzu/EXj9AZq7KhUpQEDywz
CI/8gVZT37+vt7AqiegTX9cKD8z7scY0ldvnJ8okQJMib5fKCn5ww69WCeOpJYaXk4dfegtPvecc
1v1nLWalNV2n/wIvMPf/Uk2kgdtFC8wP/RJ6RgUgQe8lan27qdoqS4v5HQ9FCst9qRMaf6ia3LdV
fxgKCmllCaSFaCjc6Sv4Aig7zdiHRCAcB3P3HcOZDhOERQfcCS7v+DWru0dOnLlqHf8Vu0TjV8im
cb/1loPnvl2/K1e/oK5nhOa1qiqhJlVLVdSaMDvnA+OUHPKro9r0QfIre12pxvZtcmfR1F0X8i/j
S3IFWHod1F17suV8i0DjPodtBeRaqW60fLo8ZtsPpamTSWNINf0dSHey0UOrdDuk4e0p4EMc4/e+
/2BkytZxVQAdVc2kaauesFMRKsTMbaVDE8HZlvzdId5uy2x1Rxm3Rl4QAE4GZsM51Jfrl7jotR2i
O0lrWWMlPIN4H0PUDKozhv7YCcCiE5GR+mTo0XLMsRKERzpXvwASNRonQTx54Y6FypccTdSu5Mly
fIhD/vwxEwc7EcP6G+XVdzapqspgo3PXqSHgwI64di9ONKjdFl+bJYMtLXo/mR+AzU1fr28j5sVr
FsiCiDSL4F6KBc9zZLRPVGn3YQNd6DW2O7UeN+KEY1sLKXiWqRFMcbkHcPOieXh7PA6lGDe4x+QK
RSCgzCBI6uqQ1iBC5uwygUqUP48Sy6yWZMRHpd/fDmXDF+SJKxoEmsUfdE6b39D0ondoKn6ktSLx
3gCwHSTjJdywBUhKei5LKvX3gN/5ees3EuuEE4ScAbk1bEARb3AzByVfR5PAFSdhsFok2Oy65A9U
HmjCErglunlfM5VLXoyW+1/nI3C5jm/lN6LqjrRVVMuwlJMpibJGGRmYXM+Y2SR9mCEYZVLYmYU5
TxD/Dp+WcI6FRbYSpeJLkdehKGblyXe7LqhBdwIZ3SNGFqX3aT6YxLpbVQm24ovDkjhlKN8N2YBh
jpkG1zWnWYqtzkcDh2a6q3bfjHTLv608jt7JdUWDuKgplq0PwH01ukE/gQ/oBit+pR4EHR21oBJW
eNJ2jsL+j+VVtQ+L0kgZ5Pm5JGE9egQbpkIjUo4CzuVEp4Akk5Lz2Jg0cQxfiY3Qb5ggox31EBom
xYt5FRsYTdQl6HLkpBzbLiqBr+29SzsG2gRFUNsGH+sDIlOD80fZOeHoAH683hTNwrHJroQGDjIM
pCtjxuT8FGJPzuukVWbifX55vEYjyHOXbhqBxQ4nDTMmEGBpvVItCOEQ+CgrsmtrcTru9HwuccOZ
MIavBsi8etRlLSlzk34GzTQ9YWjcPTdO7I75ngTcipgaaccI4w7Uai2VB/l2ANyHqfAa3Bg/o4bC
ks7klCjjO36eOby2VY36Kofu7tI4/1aq/uRW5Q9PH72o95bv+vJZRM0uqGqfGoHMzbSDuB2s51tU
EOurcmx+bhMaykr39GQWUgwXzKUwTFNq7BARIt9J72OSOW+k5OifeJCVVELk2OaAn4GhWVpCXYqh
BRirCBRuSDNJ59jMqFbDHhkgHIS9eLb2JClUwt2uT2w7A0YgdiPoOlZ+97e43Xd3mYnIHBJTMTts
2uMAfvvbqaIpHd/XX5/vh0ltW4msgiFyvx8Mjt9B7ru1Vs7B8JhCl49dVg9SA6/0A6KNN4iTpVRN
L08BRIP4RbfeF9FQ0KJiMEdsbhU7qDrRVqcJz7vJrZ/xpi95zvrfGhB+nRhYjx2DGd767/Gfycj4
prTkwtmrsWmopuj3KVxQyI7RZvBXANT4FZI/KGqrhfmwk+0/G3MfSM2PLtSwk8uvjc3DUvyywBUg
CRC6S+L4066PVTBAnki12jHI8gThn77HwUwe6GbY0aUxkIidEB3p1hmfiZEnWQPW/fPD3hO2UZHO
S5P7N6YnZgOdRvXle8u/+Bb7oW7XyVWNzwBp77jjob35yTh3rpHZWAqE5ESYvuYvaYhF6Slj+7Az
GBaAJrwlD5S6del4bQxBnRmU44RPbQcEdKrf1fY51m1C8BUdW3H5kk2wKmj50dwMrMl4WP/7rdFK
3w67G4Dac/ZB4Wq2VilJ1fLU8qmikLdYgFz+krUrXapTJ/QKaXCcUtiSIeNAiAxsuA1UCj12JJy8
zkgaKM2wItyFcQ+S0yxOSFDZtKupN93ZWk1mPq1vG94rb75cQ+/itt2XQREFGtPpznhKMhkONz7a
6iEFvjVlsSpRkc1WIE+M+dMJWizGj6OQ3+dNv2BB1oTZDmx2i9JMZZRmAMsFGWJCWLPMobA2SWUF
+oy6attLpLyzNBJDOxWfolDXpiFS+IW2lTLDWmwQcTKjpzXwykOAe07GmK8Sh4GGCR5z3Y33w7fe
zJWd644p5ypxtTGmQ1iWee/bgszMsScuuHe/0MifuZifopT2sA0SUveAcrtc2m+/E5obr8EDvzcQ
2xz93vD3+cVcSCSIrD799wtMJg+/Uc3q7F4bic7jhXCNlll9sboTP/Db9t+KSRThtPDVB2CbX6Jl
A55n3BDOKi20/FA0hjaSWl2q1mYi+5ugkA3vjKtMITt7jgkRah9RtswCjvfdATA2wTwRdj0b2kp4
eKS3nMKgdQK0DTOVtBHGv8dTwqres4FqH51t9NDiyDArR05H0SOlncQeyObLl2RIJxp7BpbunR8u
Wly2EZ6rmkhtgr1wqWPOO7D6eVzrQAVoOYvzsTffC8I18TbhN8mHWkoVT8a2hKxwfR/0iXPyR3f4
7t2yIdTePv6ICz83+DqDW8A0/u0cC/N0Ti35exTH32YfAptUv82QBAB12aGkevZsJO1jFZm+0LIV
2QmDCna4HTmrfhXcBHilicpUmGW7CBLrsE1CibY/t89ycA8zKyUcGQPXMajQUPmhH1ondj8aMlsd
/ZKqQiXnDtlxphoYOzo0iW8zSAMAsgDw9Gh1Z3HJCG0O+RY/1kOnojRwOZDes6pKP8o5mxZqCHw0
iQyBCKZodP+H8tCysyE9Rj4aRtPpLCvbhBgULF3Z6eHzg+eX7e4h24x8mcdyMB/K8+kumSMtjRct
iipHZ78AM4Hu6UY97EvsHQPkEhBj1yptBGZt52m/AYgp6pDxr4aewpp6RU/hgE+rGoksUufx71O4
aBhE3+/d+wwSGIFoKx2o57nNjVkWH5gVSMWxPEmcJbHW9kXF8gbq8luYw1E6sgT9rFk/D5NiZQRT
rAwSzs2P1EEA/IMo21RERIm61gWI74685co/EBrXBzHyt48pqnAsrOZkKRXsBjTXBTlB7+omX99n
80LCZ+vYNymjiZaPNFTeeQht0bSaG1Lj0bwRrXULs8bezWmOOIUc91LmC6QZ3bm1qR4rKDXfYCLp
hlcbOooMXZ/8jgJuAKouMH+Sd6tbgYPNJ4yGyegg4Vu27aExlvGZ5ieGEaG0Z1i2pM5o07SsVy1g
KhsRasKU1lAi9wMxlRf5sqBCmIVvY9kdS0UweBDPl3d4SpkEUXm1GkLn4GWDQZGponHjn3IomAn4
rm0poQxiL76dFvl8QoGlaD2LzjJYjOi7wRmRE1+emK8I+Wie1dFf79/bskjrqSZbBdGUuDyDWCIF
usq9qbsZe2iqQugy3d+Ti69JbutEubJIUElApp5qH6VOigCSs+uCe9/3YENudY2CySHQ4ZLMvPbG
zPxTCEQShdBjiqDfelTUnpBUsezafTL9/n7Yp7OmoJsHXBErnKm7KhgsF+XcZwaggBounKXdPxZw
/aNimcWCO7xkj/MDr8DkCzXO7XE9EFG3T5hy3By535ezS3juqqnZ/Dmb9M8/Se12si9tJiCPp4p7
CBdO2ATLR66p3gCN2sozragBCI+lIkBtJJpHT6ST/TkS0rfrxt+xX6WBpJO7Szhwfe7oDGaTzIie
TR9/kh7vZh5fRZ3bxJArrMkgpypw3DLdtKcEF14uU+ZiBEfjaN5XDS2tO0m2SF+iD5cFwrgZCpwc
wriJ09RUnrSDaStwmoxosQmDBbIR35uSmB8o3dOM+iHh2qGnmyySR+y+O20+NFr/s9uyGSODTTLY
C7ql6C0Ff8mghqDwIssLLKu6B4I7KsjEqGZHbXuYwdIUODnQOruN4idUJRNKvAQy7CiuleBOVDzc
9naruN2yp1EMVrdba57cg73pxEuEQWNBVFU4i/Vs1sjTYH70aTmqWItgUgDHscWf8juTTcRORVvt
YiyxzGRJFGb5bydVRIXrmvTdt/mW9L5ujWgysWkevYiZ55Q9cK7gyhswFjYFHIyANPyeIbTjnmnO
n35wPAr6s/rD/fFgW0f/kx/MaUM0a/o+p1Icj2DRQKRyuQI5FZ3LiF5RvMue9RQ5DRCVPJ+lXHx3
9CfbCntCVCdCd07T1cKykgR8+wU+kP8OKASF6lGh/zyVYDVnmxDiLWuFrswrrKZM9Ve2vC8+9/M2
2+YX3FSrpLdUCBauaWeSQutmx/rX6RkP93E1N/3i2KrUUUkvybLa8YIf/IQN4g2tvjS1eT1Ikol1
2gHZ7RyXElEbjaH8XjBuWqeZFA4FcFLmjjsMcPvAcRo8lDD7Oic69j4SGsS0ezQ0Y5+fXAvagZmK
2TR5UO/wEO/u+yC1HvXMNPrDiXjuMF2NxsWWzNJ9utboXKUw2lNUXUr0B9GoavUUnW6rpmw3/CyF
Fmo7U/9CRl2cIBHwpxo/3utUoFmlv+eCGR7ZWcHfglOAJHfyhzBVfte4mVQfm3kh7dyFGTi4NqNV
kYqvgfMnsxr7q6BBNMmkliliA1Uut3XbqltLjFWngHyL+we+xz4A90SlDDkvcxwNqGA/JvWD9tfV
wYBGjGI9knD/SEOl7SGJ7HqG91V7gLwxNynEyPGxJ+tlltAVxGKZl+TdJJDQtvzG5PBIHab/SoZn
OkqdkdZtbrjqyE6T6Y7XCsRpnw1qDjUvZGYpHzoi8eO/0OUSIUCnjc5XjS9R6R1oRkMgaoGHOxom
IR5+Px87p8Bk8lBvR6vuMrJNEhMz/99Q/L194P0WadnZ4iBpR4cJFy/cvYXU0iKFmI+x51gy/rpw
RwbxNEItw4eQ4xMUEFhiYfCzMs4Wlni4LnuWpN8gq/u1yQnOGL00s680lD762kDbu3h/lwLE7ofG
xXULCILreDqfBtMFCxEi17FGal1cVdx/uGV2I1SaZdyjH6uvJBMOvptxUYvwM3ZMyutbnkt79l21
XjRxyUPrI4o/8Wp4HvDnOtuo1aJUMx8+9NYgIZ9YOl4TiyP3Q1PN4fkcOTANnfL7A0fvSOLc2xsh
VOVrMuhdcdgCLo7Sh6WSMNsd5PM+qjH3R/DKEJsAdg5bcqI26i+upN8C6qP7vvzJEULQVOuQKLBQ
lIXN0efUs8FcVB/YRvRc0h9raJhHUunGy1wndkvwi1M8YkWwU9FdQ2QzJZOcYUsnSnwEyWRF5OxT
4XswqJ4FXuRl1ld9z6Kb7Y12GY84RB7dDjKbcK6aJBX3u5x82JNzDYHayKBHSZoMUqY5BXKrsF6t
WvQGm813gUUrt4YS+dM/2px7VEwTqM7JKOOjoWKNP9sqWbJqCw8gW2+iNzIUG7Io5NPonRHGMLgf
dwRg3n1sg+Mf0LdxdLuyu79L8yr66m/tBc760DCON3JQDJsitoTQeJVQ66uDf9WpbZ2fXjpJA5nG
RXN7m3Jea/rLExKymKU1V98BgcGFbCGgNqjb3qvFNWxMpsONrQ2nrq1vtDbIZAWsAVik4Zk4kdos
IbqYvujgNWPhhaBXuMiA63LKKVzvMb1h76hw5tIX7irOu/xKi0y1MfW8QwHydsYjLC/zNHJ7CEXV
q8TOCoHYa/eSjo3O3Ui7c7JbEcHI5n0yRNqflT8R0XxBUEIUt5pL0ylsWhdg0ewsZqkArsIpeMCG
NJqP3KQL645bzi5U9z9iH5cXvkwAZRBA/rNT/W7d3kyBJGe76tvmn/o1olR2Q5myBLkpAz3p1v0R
yrJ7p8w8KtypUBtTWWWhuZHcwHqbHC0cwj10Y3yqqp1S/pL4Edkz7g2tsq82zcZCKwQe6vMG/f8h
9dYUx8hAGViMVnJ4E7RSAfzaWVBm5mSVdpkz5zvGfmZvjTByPMFL41LpFIoshRtIc0bga1E4Uln1
bskCBRiSgG7k7+w8W+aeO9wdX/jsgaOFXhjagUDJu8Mup0/Wc+qXumkh2yU5IkJECw7htwvQpYz+
x+3RHkcNlyENeOWfCqkNgVbx71Og7aURV/Feamlc+ZiITRF98qX/wWDamJXLPjmoAB21bFqaspTW
txCyLP3azINTI4H7pAY8s71anHccthIOZqjmq6JNLyBWG6emYq2xoZj8YZi3S53pL077e7A2sNAX
M/h6nM8gezPisG+Shumt3yMpK2DkqHPav9KuhGAXYZgQYnP3ZKVmdQ3pQli37wEhinmKDz6OvybT
VAw5NQyTMUOXpVRv0/WxBeWEXS469IzX8IZciwg1Wauul94OemmOrCnEbppWpmSYv4b1RDSBnwyK
mFCs3Jgk1XOA1aoxCeosj/nWFBu9WpvGVd/+GXZetZ+UnnrCvA1IUee/4ggQCXkv8PmQpkgiyWBI
yBiJBGpOKhFdIzHHI1r6wkGxYYuD+/wX+cp6FCY8VZoSF7O6AZNvJIi8onFyonKjPoFgiHIY9suY
XU+uxAWsYmWAWF6g8K057kdAhXxnICgfJL+b/poRlCMDQOC36rEBBq6Vac70oxR8G6tgDoAImrRz
dDUyZu+F13lHIOPX64wuinLXATiFcxziAHOpu0TftiCYrBV3O5+1O3dCS/yAKBrdfctcMUkGcqVK
moE2x1wQbuvuiiRp6I0MW4yplNAJvP/UB8VcYXlm8UedhYZkkz71EpSqThccUxm7mt9pUly9GTxT
CHcCX527XV+Dj9zemGGCkNRtSlWhRuPMaKbfXzFYJ2JgWV8NDxT4nKvpvVbfxjWV22zuaYswrDDD
ziElN/jQP8nTd0waVkh4G4eeqSgIdOFtgl4DsrPlPdVF6AJCwS59u7H9gORZx8R5OyXemqexrDnM
YpUEgdU8ojeHvaRGDJ1GvyLRko8CmF4xtFHvV2n37Nmfza0Bgbe6FZgCCvyTErPQoOxmn5/cxe9y
8hBy26OGYMbEMFso+zCo2Yv7UUYtrfXiUFRBYwnWDWkdL1RaHsbdY55ojesbJHGIP9RvHLnC1prR
hQ52ST03a/y8Ja1HLbhj1eUNLODRB5SQVUZGeZPoY37D9RWKGWO5mreV81yxnWNmM8dlBOiv0VIl
EhBpxGGHUs53mvvU+xt1z5Fv0PNZctMNiVngRpyS8OXYfJKwtC/8h3/SpViqgbrFXfxrplMOdyhp
OqjsAqgzUERQkt+x9cwBwoF1B8LZLQ/a35Z1hrQQ8gxC6fNZCvEZ0v0kezxLQYMJqIJS+7+mcgX2
BJ/u9GAvjFNsqbRTjvKt6/N6ln12fOtrqRJBgLn8FqBuMNbJkhP50IgtTJFHlmGHL8Z0Mnsq7/tg
RgcCLiuJIk9/MjEVOaxSpbwpuzsOwaNwDJWxa8bs6pA4wt6L4pFw6UetiZlo7rR/GypHPmWx+Yes
NUT09eN9j5lfBqxN+MppyAyvdSudQe4JU1D5vjG+go2PPa3tcCfvllDMZHSVPL/waF/NJjW3CKzt
puPenDOpvXqCa7m1t4SkkxW12D/1afcV5fEiWNWlAzJb8AEq8E8f9C/scQ77eAdGa3OqnsZWWU/m
qWWVUtLG0kuToM+1MjUUqNDXm0xj4pq9qyjbNM36SHSS3RzEgzTGG/9yVSIPCZfB4UWDZ/Ybxk7M
P3P4XVLs956DG3Qc1GNlAE+kaw7qZufm4rLyi8Ah2YdiftLcho5izVadMwMjauvwvKVFs6jbIX7b
bd1ZfbKT+DbB7W7E5wazdEk+xL4ZNVh4O3mOb7GHKvdhIuPtLAwfTJ/xlWiYeStAfZMovOmgEngO
2+XrYbZQBk9UvjMssLDkrYMTHeqvIJQkP+HShlkMxTA1HsNuYntY/HiszkyAx7BNdvs5cuNd9Fbj
jirMsQ2x/bll1R35FoUYDEi8Avn2DUS5xJc8lcqpW35NOdrT7vVLviyq05DEQ79TeUBkZlC2k9T/
Z9I7qK+JB6Rzf50pZMyjaIzp49WoqDqU4cRWSlTN1X5zHsqkf8z47qs6jfxfPmfwDiMMM7w7z3I0
Zt3Rvvym6zU4jqhK44hEMj/lXm+GUJxR2C5jj4lMAEQU+59u5meiKOQsOHjTvDbpIQafaCN+dIbs
02O7USlCzkPPYDi4BCk4RZhNxQNES7JkesaIXgX0vnLhwlw2QDYv2QSWSLSDdK26oXxUFgQYT4qj
nqbypE9PHeppMfmf+Fclon0hbudUUU16/fThGW8LO+8NDADAxw8B1UuPnydzAkHvlZtr0AwoSDhQ
dwgYzHukLqoq4Iu+zmS5tEkRy7dcgTibZo2NxzJm0dmmuRqyGli9BnbTQ0x9h2d21udc1j47JGAP
i1zxHudKkh3pFeeI0IBba02lvHxOn/Dn3XJI0E/a2w297WIEyXbMk110ns2Fh0z6R5kFYhlaFItu
KJXQ1S9iJueSPVrrW3La+7soDGVGbJy+sV3ruDKh5L7Qiiny7qJ5dGwHcqDjkMJWlpTSgwppUfhh
Zd7PzFNNllJ13E2QpC3S4MvlyspJguGBSZCV5ZzSKf2RsMHkAXvPjLXQ06kY7fhMJBxAwqN7yk8I
7z/MyztHuZISMkAz9RkeTlZ1D32wLAaloNZgZMV+noNDDjeDuUwqLyViz7OKItLbwP+48NE2s6E1
VIdXyHYRNx7Txl21UG2TCrpBGV5vXFZp3L0CwbATeN55M8v19LZIs3ddaA9+Ymj8Pn0l3GDh1zx2
AAlFL+URwkcmqIo+cGd2spuG9xf8PjByb0yxygKOA2cP2zx37PWb7UwR3Ye2DpoWhJNRumiPSPMF
m47BonzuEaj/cLJFds6XCmZuQpKl1HCCXZHTYx8mszTJr0VnNe6CfmsL+rcz9gLg8IKDrAOhXNSL
Y2sgDgImnaFIvwWzVGz2GJk1m9YQgUktRcsbxvrgZDykDf0FEOAdk69+TdtY6deQ/DLjSiWmqiU1
cIC3TedW2gHuveUxcBckvdzp/hZNHgS4Dje7d8m6yQ6eIUdVN4HP+F1hxoRY4QuYKYiGLg2N7IgF
qJKtSvx2G6XMsTMp8Iy35/WGd7YmNGiZU81NR+dG2enAj+gZNyxtY7e3Qiyidz0fUF+LxpM6OV7n
yl+3jGQ5omuCDeNC3fUY9ctNokZ4Dl3CnFFHxTQ+eG5XYdCFEPId/FAgM0+W1wAqUMyp+gd3Lp+1
W3kUbSBAq11wOz8H4ZsJ4RF/FGbCQWRsxHZdPWLl9h2FP+Kcggp+IKbDJZ9tIkT8fqukmqzXIGm4
FrJeTjnH3YnVkdgOGn0uCzmI0f9p7ev6iiC1RdRPahQrSGNpTsq/1lESnyvOlz0KJr9Mhvi0AUng
KvsmRE4HMUdE1wdSnx4yQTtmKdDT3gTUOgX5cauZO+1XpS/v4oD0ISyS1Ghvk6A6FTJefBtDeD0I
gs1WMTVajdOSdw7CaUuCcTglQnKaYuAnRdsaNYJ2w3NUO94wgTP4ewjwLSsqEEGJiSaQIiDoeMMG
KFkDeLFfwOIG9i+MSdbYg1McWxV0HUrY6R4XdnubMlbBbuKl3Q4BokYbOEm6F4nVQa9/Hw1UuQZL
uzYTbB7M6d6IqjV3dpx0Rw9t1aeOaWTgu8DNOkXjCBhP1Sa+ftbxFGCAKKNoujN4P/Nt1g/5PD9a
sYYtJzdPWPsLqqjjwiwFg+KJPdzHqAJR06bE+sAcI8mQnxQPzpe0L5VPzXZPrvBbhL2QINpumkKJ
vF0em6iS1VDoP5miBSYNJL1UyygvTi3MGIwJhct119aPttrFoeMLDLIDFd0I+n3gYbLNdUxiSLit
y/tRhYdioZkmvC7jUPNvLeywvSWhkKTCCz515ml8Kv0jWC8/5L3BHcShIDI20QIE6PZZVqF/ZoSr
a6QV+CPr71HiuwOIitqagE2Pfr9tPHvEGqvECoIfJCtxFvPbL0ZO7sKXV8dTlyV87CBMnh1OibO6
0cmrIiYXyvnlCPEMCMmXeAeturBkEDm+pss88xbeTdzcw2EFvTjIzz8oYRp4+V78vtytl8OMo1iX
EamNnW6gvAroyUXubHTUkjV3LtPpE+hZ3gTp+1BvKLd0r9L+rxd+Eb9VVDk3InfNMabWW5JEoa8Y
fJLjVBBzyjnMkK6BaG1zAM6h/q4FcJqYGBy09qtSeVGj87jsPF1irl9zhN1FPHUq85/9alfBEbh2
qPXkPpAccYo3Mzqb+2nf82JbCDjnEdUwKRMyYcsd8BucQEYZfa1agw6yhJo1kyWmkkYvfaOCuZco
/HltWY3pWednC5/uUiGT+iBULtvzMl7VDnKLCmBZxUy06kKbo7WU+2o24XSauK3+KBhFgUwiy6Pb
rfcvtXteAYsrU+Jt8a4caim6MwZPe227eY9DdOfmVp6QnpAJA0Wi2e3xz4aHZq3Vl7TimofRcYXt
vqbNGLNupmXlrYsaxK3sFbHdac9O2jZsxdcls8xQwYZNTNNXWmZO0vhknPMLfGb5qmbRRmBrCw90
Mq+/JiLPKrmQ8xKlK5xAFYnb9E7TlFFaKrCY8LkQcD+UjIe52yzkUYejErWJft42eXHLDHeqTYmu
RBQE5G+uRfOIJv0qqnGOD4i7Kdry948ySp0sVPYkj0MoGm3kFpsZ6/8UsX/zwlW1xTDtL7xcFvDH
7p0q1CDxGy6NTZnVFr5bkC2S3xgUqKEPQcEwC7c7hdJk2dd4pU6idcGut6hpFxDDnIcrPK2poGXN
XuV4VusDw0VzCKWbSTbwiQIsboenxCudclGke1Xd1RxnM7btuLGnUpABFPU70iBkmrV8kQHtbID3
xdqJu3ZTGENCja1Yl6JzR1nZ6JVcle5KbYUWfU7GHoOqeNqs4/wy558+kfD6mW3bfNP+sXeOEGN1
igQ1q/mwkor7hlqdZJH+Mb76w4g/4YYT91K19iYDFAGtFxSjrpOemycm5wcizU0djd5FYd9MtlDv
vAHWhxootTN350ySmieeew7cpoqZNMaF54jR2s4+Vgvus5bIayMcuPVBOuFLfud7twlZKQP4duSv
JqCkMz3f7IOhThcqPfKkLcNr6i9wEswyXplpkklO2nBrCYR9GhbrNdfCv/vuEMkLSpLP4DbSsgpP
nOaqjQ091UV60qO9i+YaTUGxl48ZbUJien4Wv8ZR3NjNAcd75AX6c8tfNcTj1N5se/Ni5ZDwyNMv
OM1eaEF+LutGXfZp/2pXAKm8su8+Cb58O9BHUIrRhQ0HkDhuGLKcBpbqL+6/zjfL3n+OjhcID6MD
fU5XiCqvjecHgijSg1BCI+z+Qzy8ZNNSpuoEwd8dKL/sKbQVQzPmfq+1tY838a0N+SKdhsxnPzXe
93yxnGimsFwx2MVp3kBenaKIEy9qfArqEToudFbRkIdmhtXQaOD1AfWXbagOuB0vF7LMFYBFzXtU
yXwTD/NtJg1560eZvYMghV6NWVILuNB1gQavMFdef7dS2SqbRxpB7/t/x1BADw+0FZMUvmxZb4Ns
/8bsgrg0zLoJYdEeQPhhnL+CERD1EFXvkJVUYHqAal0mH80pZOoqNuYMmZcoGiEEGdDRuFYno1lL
PbTXamR0G1sRVsl2GxLIKIgUhG+oYiX4W84iG89Hn2FGCHCBrlClkQgu1Hp7fNUqzbjbEg19nn6H
EUWzSMDjUsKv0dZXkD4YGqYIWx0LD4EbG1zGhRv6ZM3qjS1VhTJ5lO6laVeZNlMGmNEvf1ogTRFq
kfZPc6zPVQDA1TC/kG2Sq74yVj9BkaLgPImkSIsJEL/YYbZaKK2PbmF+7wo8iCJHSFlsUJPhE9iI
YE61h327sm8hofEZqrd9SHQVSsWI3/Dyy4dHQpa++zGeZtIura1ssv9z4Dl8bTxOCVhvfm1bmbMb
d0us6ej/jnm003CKW3s33ohi48XnGpXK6tHYRVVoQ/p2k8ZXzOYdSdtP8Z69FvXIRPKXbu/iLaGY
BHWcJGULz12mWtkmlbSBCf6PgUirGWdmKT39bWIdb+gKrMjDdiZOzd5tkMag/3mg0zVJrKswYa66
KkM7/vqe+8BVPs0LZS/jAtGGb2kK9e+30i1A2HqLMv5WKoEi7PSxfIz4ohtEXTZaHDtSTFA03mgs
yJRus9cc2SheQh6uIh3RUMMcaxAVcynBicOlrWNzy+1Hr3wLmkrUIHIVYsVJHGn37dztyTS9hRIv
YM+yoIXkCV0eeq3w+nRvDr6mOIkT4J7YIhDB0ru3kVjS/lBzZwcSfKZ6QtOqhHZpq8RDP70dRPBg
V9tzVxm5OT2wv274uO/p+ES0sHr7zL4XPzJAdNGMA8iyE9DdZzIM1Rj4mpj7mcvqYX8UO9NzRuF/
2sNK6gcG9mlJAdvv9qgY9dtwMoRUZ11gq2c8XCqNOie15273tebb76pELosc0Pvy67ghzeMP9R0X
U7MMvERlEWjn0l1xeP6yGsC2LKCyJdUJ3zmB+3y3qJZao6C3WBnuGCVbuQ+39gsWvwCj/XtGBA+U
v0sD7I2dsZPIS8Shv7bTMHfqls/iV6Z9eetYlIDtv4sQwdQq4aoIfDBSFxnNNf+m0NZK794JfYZN
uu4tOqbkKRA1TSbT+jzsKuHkkBhDTL6h0AWQvyQXOJyjabj0Y8ewDSqMQQovOJriSywWwPbvlJw0
BwgR27kQL791+V2rIH1UEm6BcqngNeuKs2C3t6NPUVzZmpkfC190PtWwwqhVi99nPnH51TE2IIrG
nHI33kMvtamBzq8WXmEaNUKcFpL46v4fyLX+j9oeDI8fjuJ0kRtQ3GNNqElVK71272Ki8FeCQdhl
EGYTOpB8hgKsoo3yAz2pI1po+oDh6IqMlyTVo5iipB84c04RAG+Txq5TD11nZQmFZwnCh8C8tZx5
eX+MwS5AJH0Ip5xdHQeBxnz1xcFfjdVUhFkbiNWzARSr/5LtxmS6uXocZMeFYbrtcauaUzILHlcx
8BoERZHMHGtpD4T+h6QIhkv+7DS5ABTJZrOiNBJaz14ZXJSeMwABrCvFYfzj0d8K5SCOsU+ho4ro
UzQKKOP5N6igiYdv/fHoDxHcUWyKIsDRqY83HiJzgtNw5s7idYNAnA0PiN0EHR4FXSr0qOAZHcQk
o7/1e4POCUK8AsAi8HFaFSCy/RbZcAUTldUTzIVJ4/GupndVBJVga8fqRFa8U7HSVLk9cElEG/08
ug3rfE08LPJ0jFRReME/Hp9BLX/RA2apkoza0BHZX36fmDVaiJvU9QN/9gEdg0n5FFyitoBl7068
lLvcA6H+siJGWnjjLZOFlIjeoaBDxMtf0yz7pIfmorJqioc1GhJsvNGIv6JWNPcPyCWK39c78DLn
Oa1BEl2q+PbbzqwRM4V+JKMkr4d0+x74MNwSLgpaqsg9TmX3WFsC/UIEn/Jtq6AIkyRbkGGgnSRU
xCAWDXFn+1E+BR6vRwTU4eofmKvT9+2oDMuKa3uipgfP2R1JBeIqkkBanVjJu3SAUKz3BeD0jUmC
rM2xJdQrIeskGoY+LdHLur9niqkj+HuyLpDaCWMLQO0mN6Q9VaL3nw1f7RraLwUh3oDGNuJek6eh
eFFDEya49QMksQTCXojPbnLZQPr76Xy3NfkBUDlb4iX+UXPZywUacncb/8CY9qJmcRyxPA3+KGWs
QnoluFgQmGdxiLeBlMe09k7FN0Y/0EGaZs1iusCUJHnVWdZt8TyoIY1ZVO2jFANh2sSk6Rlow8vo
dkDLW7hp2yH3SGbJl6Tkqdf+nG5uK24n9EMVO1JovUrFtBagD4ck6JcgB2tOs46Jtmqy2Yf/32Td
5xvLW0wzRhwz9gSfFeluvNwfQgiQsg41I+t/MrS1YvVrOh6sB6Ux5rKEaIf3VtKwNurw019Fifxw
pOGsuunGHgK09ZO1xtA7eTqdZ0AHrjokk0tfEI4DbdG2d/DcPG7TWVxkGTAwitQb891KFD5Wl3NE
a9aSCnTGdR9iQx3fU3Q8yBv7t5a27eRKTdaUEyyVdg+/6/Y4tb6u75+d61hL1V5MM0f62kI2/Zxq
+JwUDhRm9LGCFXPHBjbYZjiNdrVy/JDs03onKRasFHWQ0UXTgWRvUnshBWFJdoeHhpNYS3bmKaMT
imyR8LHOLX+qK5MRfBfT1prwicuS5/2fa9FXh12zbwHyHsyCMAVsFW14VNgj4BhGDFh2qoDZ+0Lm
BGcR2hWOz5jEDZ/pTyF5U0TgYt7qsLiBNPzhcTAtLsieFdS+K6A7EBd+4gFVtxe6C41aTGqEDS45
nTU++tNvVJ4eNEymyCF4kXOsDjhaih0vWbe/RO9owy9h0/5w9iyOdhJ2qDf4eIhLTJ9t1kMnBlQr
mpu/IUWtOIZ0NWUErxPEmWzJoGy8CElbOBDxiOvmbQKz8TrMr8eG1hxS/sncVDLl04uj4tHHM1VS
j6y9vgibhfNFBXPQkpweCjSd95A/OBdeTJvQKmhg4YS4hWFNO0QQD16r/sYBcNqLwLfdsRE+1sy/
O4KPfSwFdTp+jUxhj1nUzU4IuxKOGCzRwgJhmWQhf32/kB5ansY2KB4n222jpCELtBDZQ6XxAWGd
SWrgqJq9LkCwsyVrs4t6UMgGICuR6xS6/wOFDix3ugpS8I5MDqXjFtwRpyKwHiT/PWTlhqPvQtal
EiU81zsXeS3LyNy4CWqqKnyof0tEFF5qDFELIG3u4csQyMxLizKiAs8uDr95lzroal7r1sh7l//0
RjC+Uk9pAviwsTt2a1JFAWM2AdFPsyBDoeWcHpGvypYcTagPZpQxsvLJ42oyHeyGanFzSwV+EA6F
sOaL5e/PvrFd4lrLjiK132zjTJdTIEBMe5ssLtNuIJM/KzLRp0jebJIdvFZYPxwvdfdG/GqZV+v+
doqHvJxWhO7EKJLGOjSMihXpBRKR/GD1/lsAQSBYe/Ombx5f+k5VLklBrREjGlpovcgiZKBUVm4i
G5I3EaiErFH7Ow0MIHfF0FDrvD6rS3XU3JqYR9GSTG4Z/oW/YYJNcbP/zLe99XeZoTm7s7u+2WbH
dKYg9t8UWOQm596iXw4To3/HHQzVxSpBeNPQgUKo0421oXthaA9WFVohmNX/HnWt3sFXBWd77UhP
JEYukQz+wWLXMyNvrpLris8RO8U4LooyycxKkYJVPbqD2AOu0acn54YWzGqooq43chKBPpU7ypHt
29bQGCO1ZCm6qzLhgzZu/rwlt55F6n62xpNWfIq2d+7+ln3UWDCODpl8hPDAotbWnOzcx9ZTdjOZ
Mi2X2G6/LvAecMmHTeIDCjXWsWZIGY+7kjFJVB8VRPsxzccON2AhtDsILUCDTLE45BpUde0bIbj4
daz+L7q2fk66TQHdvorDUuFWhzLYsChYgQKR0cPppV5/txw8n+aFKUX36xehGvv3aOJ9ZKkcChP5
tOBm2ACXurUIdxgFNf6kAk6y8q5KuzmlymesLcbYOEhemkTUUEDl+6RVM6VkeVWZlxFI0YnHXF3R
5I7phV3sAg5lAgwWBwP2wWeWqT6eo2L59q+RlQcyv3Ule4U3L7HjDkI4gfxuudBCCOem0EzBAsgp
AyYlnyAxoSeK3l7aMGyR+/tLRJXu0ueX2UbbuZmU73/pck8mLmyZpQ5OILuJN3bEfUtU7D4s6YZx
Tjvysn3MHAwj9h9+4bEm9BfOfqaFyj71uNah/aFozkQvKhuSOSigVGJu7Eqq08qsD1O7f9Aan0Et
ysiTfICNX3ASn2IKnc9eYVIUOVYdgW/bco3TMav8KpO7w8RHjGo9TJwPaCKZdgG06qbJvaUr/3I7
uJZAOYY4Afcpx9ZZtTi55eZhnxnFM6dzcx5K3iyD+AvpGoa2Bph7piYJYirqa2C9N5Z0oSm1zFoo
wTVt9owG3n4Aj2lz8FUreTlkgT6dPtss/78a/YdyI7NN/fLXzRQP/uziYcYR+8BwJMVjutRDjilu
9lVCQVcxWaW8nJW6TGF6ADabUkCVVRsEY2M1t/0aJ1jtp/XfaJvOJWw8y8BW0Q8zJDGO00VtK+/H
ECL7umpNP8HUQ4bb1pDKkqpogfU/tQrXr/7LNvplXNTHP4NR7My6H6uBB1RzkktX6GX+zh9FTAnC
FDmH4TKJ7dRVtI3/h7bV3B52cEbxp8XXBIMdsIWs9+2Ek8B6QSCM9/Ze2d03KLLuXMZg/FEutHjn
+wa19VixjYdcIY2jJcKdCh8T4qImOkzEfm5iIuqTNVYzyiHcySGPFYHYDUcHv7VSHfncGoLtDTrh
bGgQ5ws08ZT4xTjtz/d2SYkmadkZloBR05x4B4mqedaZSC030JjDgRttKMHQRiGbyCDRNCBWjRL3
z9m8pJTR8FMkVtvXVqQoAhBWmDOtj13oytKJVeTh/flrxE0JojYDJ3GP1LQS/FZ//utnEFjYoEya
1LREV5mQcH18V/DSjV3g2wD6B8PawftehUTyDJ36NNgzXua5ExsUGfYu/xCHlGJ38HRL9C9fHg9e
RkmRT5YbajN/5+5vC+Dcar0n5YHI6uf1BqxRg0XeU67e0AY2Ff5O0jDQrIFm2tv2DWPwViJUGSRn
dL4B+cAkeCEqUmT4mTIXMXc+Y/IRK8oUZWqqLTRUgwYC485ABlw+DSsUy1fQBzgUcEU+O+iAwXm8
dJYLJDAEVbvoLvWVkNoUTsIVdHUKBCT3VkyjH3Mcs7I0KS55ttGlKnFcHg5YtW2nfL1d5C56XeJU
ijDZLGJOoLQttDbHVaK/+5K5yTYhpVZTtOSWhDVEjwppQgC4BLxCyoIFHSkM6mpoYd+AEyy7N4kP
REsu5vxosLyvaeH4OY8SNPPE0Ny/5pwekf0ioLl3EdAceYfniLQDtvka/VG8jbOb8wejONUATU8F
nPC+pijhyXM3sxNqu91bU4tmHQnV4jO5Xty+J4VTd7D61QQ+tdslMH6vE7wzNyYSboiaKlPlIt8e
SSY8zcBZfgtF5lP1Y3JjX18uXlkK2+BPwyQOy0iTbDL/dZD+039x6PFdFe5kKNYncZEfzscJxonE
4nbd1kP5aLBLGqQGUwjpvg+g+x2vNU8R2ceyUoHzamEyQHpSFibldKmWlFUtu9MUr8iI89AuaD9C
pDzhx0xUtWV9t1/RdrSRndd+u5So4lR3t8BxS9CW0Zp/5qYSbGHUGS3Xr3PJtPp496XK6Oj7N43d
rk0Az2psULydY/0T0Lm9bGC248BgiF6ochKhZVt8so7RpaYDGQnjqER6H6bjGXwDCzPN+UWCFYm5
cz3LNsJDl1KadzRwQjxor4wj2RGJ8/5uEQJxhLNzLWDsjdVJqDSK0PZ/rE7sy5J2acTq1WrnfMV/
1P1DxmfAWoriF3ps+ssW0V+jiP7jfEyTk3RuXAwSiaNBSqv6LAcEr0yfZ4Hmgrf8F4wLw60EqryE
NZ9X2NAyzTvGFugMFT3mq6caGOavczpoW0tf62273oay5FFxL8ZLVqNRbcMJ2F3UHGlzF3zBITlL
bAWAdQU15Pw+e8uUmeB/N7x2HDfHpXNAB/xoCLQr/KxBgdHjhPKPmG5ftHbqS3ozWYLLyoVlThJ6
Rj4GumRnscv7bnowNw6Z+qRqY2S9yo0QjveYMnwjKuWZpEEQK38i+7FizM9HHHhfLA6Okl822B7W
zzCIdNRQL3R+0pAIhGE5aAfMpY5bZ+Fjp+K4G795CPv2hBNxD4KoimycUyG23tHgpemlyMWmcWf/
N34o0ymF1jbBtwDflA8keW7zw1M5YSKRh1lvESXEl+5KZ4X1K+y/L0Zxte6rCcUXbxsMrInLvfS0
KRlJV6Wg+3JzDiROvoaG0KxvsrBdCQhJ6psbF/U19e8a4G7AOVCv5J8CUMcz0aMZIuLlWD4eGsGZ
Q0fWEJHpUKkk696YEKLmt2dHnxzd+nQXDMZoCwAe5+7CG90LP98jrCJayDPKi9ViLPq2fS40+oeo
x08pUyHW2aisPkAZQ72A9KkaeOY7RsEtX/WTd4qolXqKLpiGznfCmlxSYzWH19/PCtz6+NMf68Mp
TsSczyYXfRcoTdsMI8ulmhkTvJj3UDZxI4OQm6kxAs1yJtC0WZag7tmDoStQTS6XCLYVHPLkPxXw
jybdYSonaNCHN61n0jvZJGbyEvaqRmZdsNTipQ6qdWQuST9Y4o5p0isS2F3ipweo3oKjvS97jQLf
lXeM0oWZYNkvW4K4uFsN34OgHf7ISYdwC4bNk6mkQjWZOP4SxGOP6gVknfV5fSGHY0uIQauPoMVt
9jCWZpfNc/aigyJX5Dc50dxlzt5uuQrF9LRbxj5oJGWQ6ReidAm1PUrUEwX49e5Lq1LG3jvTV7Ta
naQuNKCkjIz624MS7TDNiB0xKf8vaWweH9KpPs+RJfDB92URNE0SZmls4X2v/eIyQd9ZgadANWAV
KCGLZ5fIibTpkl3XP+4+vrFK+ahJ+H3pnrXnud0xNr7m4Jlfc5FwIjE00waR3NgHmUS4QcoeXsxu
6avk5sgpQbEfxxMvrukGFrAB06OsnasJXt5X0PV48CHEGc2WcuaExY4jxk1qQOwIbUsoZZvcBTtm
PwirRx4KGjarHKxPbgLClGGBT/+nOfItz6XhZXheuxugOZB1LnANzwfdadj63Y4j62X+GAPMX9IL
uDIAeNxx+ML+f/Z3BeewgEhWk9Qfe9rftUaHr4vzU4+mBjFgKzOTWtkXUX4HSf86qBWVCf1/4pw+
XRcooZO/X7OAabdDJQvh7nYG1JZZZVAAPa4P/dCvtMuPJVZjN/m/tMuHtQg60ipb1JT61+mHU8MW
pAFpML2dHWp3SQyeqlmLFgdPmc8pAKFnqM4rQ++kcjXzorPsDVjmgGvO4Fja3v02yNhFiiHSHiso
Bkc98kyFyzH5BJGVCQ4BFqt2/6d3W2eeMIROqFFA64OQDpplFRjAv0xOTDBGYXZ12NrEeVYh6GX4
DxzLiTy66UMW+rz5aqSCtnjFwLDkNEYcOqlJ9drNZTQdLOjl3cJWMKa/newNNN3vBx7i9hH3uC4+
icrez9RrG5WeZjXM5XcHbk6XI0LqtmPkHnCHYbAW/QTZ+AkCptYVrPuz5i8gbExdFaS/bB1mpUJ4
xuKstGslcXlE3tU+3kp0s0ubWnu4blCsiAuR1tmBTPgfgxo+70R8n78xqFHLaVoHAzYc9Na96Kjn
vvmnML+uDuYjJSd+6q5SrLA6oHN9r7sYsN+iz+9vZOuEMa6KMXybwbK/6bJcAMYRKtftPL43Rmq8
oU+mzGXFUWIiEeQHDJZjsJQ2WLRa8YxTw6h8i2YMuI7GNFVAb5Ns2P1J7ckGxhlCL+PkLptUqcUK
EUmngLwl2tVpveGFCZWDDNW1OH7tj/UBBVApzb9k6ExDEMd/IRZwKG928RRM6dGH8i6IVkvXNsm4
deFdUhpu+v+wwleF96E5wbdznrgh1tJkzFKc+YkARUazmcZFyJdKvvDaK13UrKdqpH2q7GxFoq7f
piQNfzzB2OnT1IZjb4zEf6QLlr1bnp+5zgGS8mCY1A3iQejlRlrJ2HLpv4jQqZvxgbv1Xd3FeFr3
lNuE/LyfJRLZwN47+UfGEE7U9GlfJ/sFpnwF4jm7cCgO/BIAApBUKxGndGTsWZuEACJsyOjCdyno
ni0Y7e6LEzdBcv9dp18C3a4CRRIGRC+8JLqnNkN+NlClU5ODDyySGF1i1w3u2uev2H+HetfrOen4
n+dFDloxo42pS2+n4Sh/VQXCJH2Qky3GLKwqVNVuz7l3aJ1EW1cSo/a/tCGeu2xspMerRA6zFgvl
Arg7w5pwEg0ZDpJX273wEITeqOTuj1nt3hra/Bo4H1cFXGh57dvkSD5iScJ+9tOLT8TtCM/90nkO
RDqX052cr7KIc4tJuLhEAaJY91tVzYtLEBV73YiNtKFAHo7RJDdlCNXhAnJcxzgGDVjnTbwuW8gG
N8wG6GyZNTA2COX+OVDMdBE13kpiZXLsPdNCHs4c44VU5HzGMIySjQEpitCv0boWCWsP/vCKfQUr
1G9Sci4t9aBjbFYer24X3jEyFjRT0lDXwyTZv2RCOjVq6yVM4lRPgWjFtdsXDLQ7vm1R6E3NA5J2
fFWo88ohey1Y8PBP8O1aI9g1APgT6cQwG1p3rjAKK3NHLEUKRB4HEt0jVTh14Ay+aahy34zR3hSM
H6M+A9/qswZvBKenPg8aIEzcvdyLOIcgTj7GwBUE6YMijLTI40I/Hw1XX71HKnuJqCOuPOrkE+zb
Ri62SRxRM7HPD3T2Xq5niKZuMOzi1dS2nricyj0QwRXOW4Xn4hiUIZjisdOoShkGpN8XoQR0voNA
TTjFj8t1EbKZCVo4dJLlTZSfE7jW8kYbl2LssA8PH2lLHQpPj6tOt7HpA+ii84c9dLkEErRhucqI
UZgnV8YzAeiioaQQH9cuFdM7JCUDacgAFGmLq8kMPwys8ck8pfCBQrqQJdHBH53nHiIkTNI4sHmn
37/N7Z8oGIM3KUEq4aU7xau4+a4+rYAaAHcXv2njZ4N/9iWXyqNAgbqFPibjHCy1w9VA0ytqUZH6
K3MfMmL6WOS4WblT0+KovX0X53lyOq17RStDzRlteTJzQOKwvcVhfcjHIO3lplSYv61FHiP3UJBj
QoB9Z7oS1Dn22YCnX3uYveS5V6Wkq1en9yRoYAsdmGzRKKgWKkI81Tf2R4Co3fKAji1DnoZDMTPP
qB1UEyFHEYmcZ1uwt+LKytGFLvQuXOVPd9t01iSs1CSzxAl+q0Vv8/Ulk7zfnmbr738fBUchRpf1
I/hAJPhPeFsjyHmXBPEl89ULytLkopelvrzr8WyuwnuQmG5pJpf2+uN4k5Ag1Rjuxz4zeOBDw1Ul
vpTLi+PFcHQZzp9CK/9HP1G7QkGj94ZDCfPGClBzliZjvNAnjKCCUZFVHryJ7RnGbI0Upf5PdLU3
uu8kOgnHl0fWTbnZpAPPdeALuK1we4y8Ry8h8RfTWClicR8sAUn9+GrxojcZLhuBuyLj/HPIwD5p
1tFgOphDf0oNAD41I8t5yrKHcZJ3wegruKIYWje45fiyKfdgxa5Cu60c5S5CBlCd9IK+yfySOUrc
XYiRTOxQHuv1fWwIiFqvvXNV3wWAHaDWmZvhXkC2NTNwyYSVVmjDHfctWO1LM3K2bdEWbygds17v
V1x3I3Ma4COwh8e+TR4eo36vm0Cxp7ik41vvZ1VFbbas3xWFHNmDIEiQ377ItoAFsaPjCcHkcr4O
7j/ujh7S95mToTq7k8Bhs8uf5gONLVlr4wf5PBdJd0EK++27huIeE46TeBZeOVjOEJwcRPJ0u2Ly
XcU0oVqFzNcz7m9d8Va4gWt32CN5wKR6pqXtVz0MbaJWaAWDMf4oyk6ASDOKR2UkfYqKaIq1OmuE
JiHdPwIcKHJrV3FUB19QqEhE7Z68B6AHpkdnR4/qdjFuJQyqxODggt7r8W0vaZBxmtxs95JN5170
catUAaKQNqa+kScDGr4BpLm0+Qqa6irfKX3mHEt0KFtFkv+2iIpgsYZsmVa6MmRn8x+qzVx/17QC
XEK9/udrPi3cGcU/K3RAixqbhSADWhb8UMsDELMklQchZ4m6NqQFz3NoOmewR5K/A/ZBhAz5547u
emMwjeMJ/8ZwZdwu76DiE7ddCZBj8XgmrW/0lPFH2FNsRL8ztVP0Vzk9sG9yiioIHvI4AjgqYUAf
WAVPB54S5C263VSFBgbc+CIRFKb47tZ9k2DFocD9WQM8p5ANrDbP31A59btvYIlMTlY15I4Is56q
B77EeiOUVa5LZAQipbDl6u/+dC5BBSMu98OIPykFIWcKdXP6Zp/BIruDWMKBNZqaaUagHjt1MJZz
K7NPsBOy//i85kcrevqMMo9ff/NG2PzrS76TXvhRV0ie2htSsWHyFvEvGafwdTJffwoHvbs952hH
xITAx+nJXg5kr9emA106eNF/nnpVHyTxREtgGkvp6awFfZqdnzIW9s3xRFav7pm28/DB80JKWMHd
WOkvw+HK/A/ZPQdalXSGQ3gDuTE9PNn8wSiWPlatYggez5BYpkJYBlD4iG2QgZZbndtUL1pC+cS1
u4LKxeB04c2WIZ8r+MUR+b5KOaMRvOhuULN+eGs3QY/egR4EB9in/9ESdrKHMIhg75vCunMvHx0f
b+wyqsH9IuNzViOYUlSSPDlAKT1VbkeaUjjsSQnu77GZ9iNLvGK1+RJ9QQaYhv5WzVltTia3xIpm
PtBvwiQj+yt8+Q7m4PmzSzNn0f44Y3hyz2LH64ILtB0yfl44J5rV+UfPs6r6LuWN4tTuTJXrEhx2
ai2qZ9XFAdKLZBJfndnCiSZ7KtteZI5T2WFLGLdeuNfV5Y1IuCI71D9mmiLYqD8bmDUxIIXuD59H
zfc+FkwyMZft1iQ7+Jj8r0zvnWjt0+Tex1XZVPEO82CChgjVhG3FWab5SHFlvjIQWTwMmB0wcD/u
/iS3UCjKd8JsV2PeJ38DtmxYs9w3SVEFiJZ2SJNosWW0/uT/GwdM5u+np6No8YpN+JrUs12pOiVx
MTkVH9450dY6DgAeCZW/fik2Mn//P3bBYfoSAXieAIVajmTP7SRFXoAy9nKp5Ac/BDyref3kPicL
WnU8jjK2XfxDnx8EKIh8MmpM2DUHO/j05S7r3XJDooK/hCS0PURD6aTq1CSsTGPWW4qrCW31V/VR
BT1qNrjFajOWHSwhu0vzbN7m2ONcuTaxJCR5/wmwa0g4sT8AOvUXLK//0VKnUa7r/KOfwML1BPpD
pbi7oVMaMcRdoj2R2m+277zMgujYkI6tOpPQFMrBzCFHsJqgEF30Kt7lwEP4OIAzrzh03LyNNQS7
HgZQ/Gj6sMo2bqsbbXjW+cDpSuN18RtdXR5Vgcw6XnZxzO5T5De5lm4JSb+RsxCDD7yd8vJXNAho
uM2gjCwuFElcD05W+QdAVuL/1yltTbKGG9joT4X/ah39N1wpATpqrvGuqUEX5YuONYcnm46dFhHr
dNiM/BNSMvDW+L8LSdUsdBXAEYkGmm0AKxxFMLI1MoMDVt+7TqQGNpH9I5hMgTRtmYK6THfESkUy
xdnCS3F37A7y2Sjyr2JRfyZd7wcxBL3eHhVb+GUu4JfKMkHzomCmeVcS95h3wArdON6XmXfAVKtR
oiMgEiIW13pih2wdfm1HMIfi524B7OesUr7brRNeZBj+WDvQKn50FF/f+OcbdBaydG1qsCOQ8B2w
exFU/dC4yB7FUAySLaiupOmY/KFlbf3B0TIUt5PNaeMNI7mqbjYPucfoewPl6DKy/HD9pRtfHDRw
Wnn0bGESJzS+ULvsyc0DPMy6h+Jd28cdcjJdWP03/R51jvgmtUbBNWIf4G27dSh3lqyOlAyPJGY7
fIemad2uhFA2X1Tt67Tquv/JO3aQa9h2FEm/TuqN5bRXNNk5VGRAaujS3StEuxRoppZ1nyJW8C6s
JLB9eylBEEcNcxfT9Bl27pVXS3taZkIg0S46sIwyyPVD9+oY4NLNGEnJaRpJ+ICo/w5G7KEZfWiU
K4m0bFmUWWid5R7ZkYzle/ksFdEHQx4cK/7CM2DtiZu4WxdmwH0SshbXZR5tR4c7dt54I++hLCEE
TzDDTRJKViffKUufs+sypqL5TsSmpJ20GqX4J3vPho8q9TUaXMgjsq0v4HNbJEhygkBR4JKt39WK
FHFSK7u9fcWUMEwptPGUV5SwE9csdHKrD+dq1WS1jmT4S6jy2+VQlXuu1cE1+A9wHKO4+XZolr1/
4Jq8wFE+5Tb9XVnYhgZQFwKGz/KM3jbGERMzxPUEBO6RqPRcoGq6ab+QjYHOtwDiheAVlJ7hUz+C
TlViB5/cijv/jKeOzIy91bzFXF5wFCrEp3i2i0SKd3P5p5a94AbhTbQWuewJwGqvWmUmTXM9Oo4J
iE23KqX8N5JjMFYFAkMDe0G084j5ieRwUK5jr2VP4/KdBc8bYyWVbKqmlzuJygqhnfZ2XTDHcN8w
ZRfcQHoAzZkF4QMWnNPQOKMvsDBUWJozznc5rD+7FVfE6Me0eD2C45HD6ElOa2MLDKhJ16/S4RB5
TUh2ZZmpKaLPGQFFcJhnfLF4tMjBwSL04iwAsdIqHmB3pEdKnpe9RqHM1oUVtJ6x9EefpB27vaIk
Ab9J5ZHOK6WOySSSixFL+sljKO1CJO6joiFGtTmXHnt5Nb9aoimzpQkOEu5dwkWO3gHkvfxMmEpZ
MWm1RDCW1NpNoBKky1c5cRb/WIxfG1sa7SEmoLi2UASxHGzFrYR8ht4dROG+a/PnukTuAmzvSZ3K
T2SHsHSJHlmhf2PRqATfI6R064zOvlJ6HBLR4ozYojlCpTvP/S6rSMDQN93pAvCicm4snj6qx88Y
VttHC6n8hrR6NNBRsDe4si5p98B5M4/PR1qz22R1Ei2Mvrpj5EAfzXq6FSTqQwzAoUDs9O3KK+ka
ZcKXArirlRzSw0PaWgRk9YAqdLnw49uW7gNTDNz03hGH3N7UhtfsG1WO28B3rvhEtVTJFr0XrmPo
SebjD8Q5fL923nsSFYjIIKzP7AVZjWHeoHdfZXkb4DKMsq4Vn9F5MYH4FwQag28jGIP7IDhBwxc6
6iMWX9JdpVOQH3/Iv/DJXyCWmaci+p+Cb6+Vj4ruzWtszdz51sT2Tx0IkOXgtjjec/ZMsFR1x/mV
s+voUT3MwVhRbq0werfuXdL0985czzYqccOcimzIRHmtWmlEGILh3DRz1QvA1IQcKmuIgUEJxxDq
GPNWtrnMHWLU/ITxrScmryo44pSkkI7z0mobvSpupjI2HRQJjOW6HChB2RzSCnlNHjPBVbNdTxN/
EnoOGWyePYKU87ZxMJfSrCvjpnCU7KMtYzzZy5HJvCbJDOqxAa/YzkGa7yHnzhDZyfv21805WE/E
48CkvBVCHQOUx3+m4TakrygKBqmPkkOeWJ7FAHwtRxh25GELS2Kazzn050HIESDoXIYlTH0Ehw+t
Ylm5zaI2kRVQ2B4V2vpfAsPAzlnvMoxSM1mDlONd9m+13gz3j+sslSPPy67NFXP9+iOj6XacaRGU
p4AxSczQ3rAC1TNCdzobvn38hdRWVgc1KiAOhLeGzk6rFYggvAkAzJItAi67EjW59JmQPucLmLp+
wGbVad7JOWHEzlABuI9CkYioKOXbni0pj9QaPeZrAFetOV2IVPBwmqOvKejC+apaXJR+wyEpmbF7
KwCmM27KT9p6hCLJNjF29jVuUwEYanSDCTOAsmz0SFceb+5coN111/aMLYAF5RyVTlpz59gBM0LN
wIoUq1dDViioGHsCZPJ6QLO1mz60Jr056qbxW8Dtwl5LuRCASTL6z4oJlEadPUdDVhQp8Tp1Ubp5
UKDoFiv6Numf1MvTRVAlNKYljEmzMv+n6Oq4Wi4OPMRqUop3NXWwRadsJsE2yWk8IOxeTQTsvLP7
zTzq0szB819BiQp6xFWOtxsnd7Mtp8YtdwtD3Dogw1J63rclmsJoF7AyztuhXI3gzaz1b93afyy1
oSif4B0tSiwNpgUZoLgdq47pLbEBKQ13XraEyWPaddFVC79kQO4d3Je0OM/Y72nbkTe00/iXtvWN
zC4wE1tujgyubdcYyqYl8n/q5H+PQegcD7AyCmsXrVU4OANlVW1xiGMgvBTKJUW66CFt+ngLmBxb
XMg6mQ54U8o1qGWRIvhx6xsZIdtFULqUG0Hrg4LhZZSFfLvXryroEbJreVXUT+g+UE6uHXzeOjGM
JnZG9yz0D/G/KOnVd1diwu1sXL+44LDHzzaU8nHqBOCtEh3N7SGokFdq/ThIklUIAO0481lJumuK
9hdeDwCGVJFwcfLWFCB7ej+MRzngRXL940dQo9K0FusRGZ5beVFTkAaFs2n/IPtvclIiht75qz41
EoKFU5bpFI+YnBtYkIRphz0xuKpnORQvdKJOXPX+0YXwpfF3SEFZ45Ullad5RjaiphXTp9kimtF5
Se8AZUKAhA98NFBSdPYsnOYi1nOAlAoFKyGHl9XGW4ncJaZi/G2vAnW0xnS2S+nVKKyT405ylUVD
lseUQzzQxoHGL73Qe2ZV3SgDjFl+H2SiE0FXcXKqq3rZoqlv5Zqy/qInuzgUyRaBXlke72kykDNz
kOq22hals+o6O/arJwtDzhqP5h/RMBdRz90n+AsgxLOy338at35E1kDX51srXigGfzYDiUcHcEbt
tV5dn0z/0PIGszoQelnKfZZ9mi4Vphv7A2HyckWyVbQLpRf52pIa2gJLrBtOsKRhC9e/UDX1CUu+
qzDxzWjqOu8FppqapQmbn4ugP8Hl5axIndOiusZfFkCkA2CtFOj5U74abCmpJ0ZwBGWCU4426FPP
hfuQIh9IsIqh8va2lGAEFu9BORbapYpI9pSggFabYzMHYa56GLq75d8vCT0eDk6RR58P0pQsFwab
iFM4NKi6reDVx62poEW5kYwyNAM6NHJqMZxF6aldH2cT5sYY8jA3hMa8PU7kIMRsXCx95XZ5E01e
QDdGvyUZ3ix+IzC1hOU+cVarHXP2r00+40DVdfeemGfXuT2mi0DyhuUACR80eJmYUGfx8S7q7qXm
l6rlF7Z9fOkEu8n6OtXVRSCmjtJHUbxSBFLHlB6bhMdnH291oGIfVXwIEdMj/Z1V5mi5fy0l+DiJ
yUqQ/UJE8UNGN696iA6LHs67wJPJBHoJvB5iXhgsMcXlUGUpVOtV2V6MwhFf9YSE9fatK1HMzw80
sje5dAUGiHlFBRkd3CHKB4XPnBsZi6ajg4s+Kib/7qLuSNtb4t/god6FE6EdJyghrS+94SUnaDci
ZsIKebTMLFvID/kzPFL+3zZRF0QykY2OkJ525vLoMxalcZEmeLXAohn1aU0/7qgneePBU4iwebVA
SczmL7efal1HJjg7u34ffPdURX7Gm6frBIMuxOBWmnwqs7GS4+mn5yqe2BzWPQuqRfxLNZC4rEf8
qx7f//LZ2aEnQrgb2YTrKnxTFSG+XDL1nPtVAzB07Ckka5t1L/0qj9h0OXo4kC3H/9bBNdd4RHPB
u3LEKX6RyiRFy57IFkfymFGVQXyk8R+jOf6K9qTDDg9AmSuiQHhhfm5u9hEWEwHgRWbmeTmUw9Mp
r5fXmxzcJPwxWZ02CW2R2gKDZV0SN6QRFcRr1+PYIXJ280a6Iud2LgKaBFGMYLzV+gvT7S4pIJj8
EzhFbqbAtNhESJzCdkHN2wUnVl8cPO7ml3LWqjc5I2kxrauN5Pudk+DbF6gMiK6K17g1PrOg4cWU
KC7lV7jX8D2K5A74rRME/6PHnbFBuso5lpsyoPVSr7+NwYiiaIv1hRVpfLIaFtZuiWaySUeJIzf5
c/NIQ6ze6XHBxJnysJbwoPKlf5MktVcywXxSoZu+pezinrptdGYF1+QEI90BJNnP14wHqvmuyyEV
yO6IYH5shc+B/2q1Zvc2QCqV1gU2WctkbV5PBX1tHem2Ml74Ub0iE8MUgnfUSg7qKaSJ3JKfzQru
Str+uOxxUMEUmB1S6Y04wHcKAw+9wjjGARDSAcmUndqzEqxIQzGROU/w1QTCNGjkI05Y38QViEYJ
cd7sN7/MTJQABbPpAtGJkaFMrhCMgVnd2sUWxfxDtzd+0Y1ELqzKL31qNJmJJdoxokKC+pnxXlEY
AwXh2Iyq6e7IN8QccQaGHiVOyAdxx7ShIqyFJML+HGwReFzk1XcgO322tjedv7o5+Z843mBBmvcu
QkvMIAJqzhAWZOFodK6+5qzdI3cwLCePfDq5yanPbGcHNBKZy/2dcnRiHj/a6jKAsZTv0Qd7tsOt
Hs0NP1/IXhuEAccSa/tu9Vzug6but+0vpS6LpU4Bf9dqyQTLwLygB8MANFw/AwdfQglhJZGndsIM
lF3xOxgwP1dhPcU8gS7+7BGG2OLGMwweyCqBS/rXBmmy4qIt2BUy+mCOw2u5tn2xMpJsrGBLCKGT
+mKuVuGaYOeQkZPYW+5UN95HjXCMIxv2FLrNcEIOBGXYNyl2qa5C1vtE4ctmm31nQCAarAi0iuPi
07aVb+O1aVfc3fipXkDw/rmrD5wDmFEjqmI4RhdgKl0veFVGlWfWhmalzxhtjFS19R63x6REeHmb
7quPer1dIhTvePIzYDPy5mwlONN1k55XPX4oOLgriT/TP7jGRmamvlDYbWUOnFKbGLBT0s38x7Tb
JZaGqzFjM0x+X6XRuH3Gf27xfoqoQHtVacVKhSCOKwgfiWEa2a4R5tVYPVXuNeTu+OjBTXZbjuOp
gvo+fCiAnL6A9g9LLsMig9WJrdZ1N5E37Y7icT84YFmLLTK8Spv0wLUAaUKz2fg57DVTZigUAe6t
qjFYVNjWpzVY2lSVwpkFUgJkAf0cNN0oSOCFSS+LT8cSQ2d+TuHZC3KCbLZoerXCpZ4UIi0zmc0S
T7FgMW0QdJm+3EkYCyoWwYUpBveB+uWjjpPBJTP0t4Wn4TY56st1uH8UbdfnprtUGiiIU8LdSRCi
MYsitEqujXf0x5xHGTMg1i3IPRTrkjt9P66inFG0fqlhvDQaTOVbvgPPpiEFUiccFQbSDV9vSQup
kiD3eeEVcS5KdEN/p3PqsWy0Xsr80xullijNt3KyefNyx+XZsCNfSBTRbLPn7PAbF79XXChcvSdZ
/fkDVMJmA7ihfP2AQVBYRseThIx19iXqcABt2o49WyTECwVSzxiXmtexagNjD8tYe1HPsWnLWUjN
gNOsNxBXs8jHp6wqSKugIKcVugEtjeK5vDBSFDHLYJqsa1Q1EHL2XVPUIMvHPg4G6iHPgC2OTldn
WVoNku5SLkks2RRd45uHyk42hY9sEccs6/freSXjNJwbGc/1jog/xav/xSTMdcWNaY1XoPomHpFv
1gwkoLHil23pFWQZU/QwHLHr3InKtLcq6GRWUe36Uu59wg8BCo6VehKl9XPxpnLGVTVEtsI48Y9g
X2jcDdWcLjq+MXAJeR0laynPYRFcC0TyuyeLwR/aUJq6vUzFpQtDSiHxFSyi1y6g3xTM6iuo1TVw
VyO2GEgeVZhu1BPQtCmyltR/edFOcnldDwPjEUFWHbd3fL5IacPfbvYWswi+wl6Ppq4DxnwXii3O
7hTEw8WRRA9NcPPkPAfX0nU4ha+uJFewo6AuGBJ0xja7fC3cGzcUBKWtxm2hQOmlzA0tLOiwISOw
JGHjqYKQ0+8zZGRURpXKy9FcrE9DBpToxmdGsyH9j8cAMCInvAyayzdZOjtA0EB6Tm1qi89UNjAJ
+bjEHlv4tgYrLPGJgmDtWTRFxizguHOOsBGP/Usmt/m66skVX7UVqGVPKki6Dp+LeyUtpOEjjHjL
Xw0oYsGKkJkJKidkLIe3BXrSla1GJ9O30IDnBH4iPGrOO9IwL6u3H78zjw7ifPiSU6nYjcHDlxTp
khp9ehz6pX7LyMB2GOy/ja48fnqrIB0iloaGbcSZ1eebGM30rC1ZhJiCAixZH7p6njj70v5NaUQ2
3EKm5I+1BlGXy8aR40jxWGY2tAZf7Q8lQOEWjoNo5+Fz0mRR5lzUuUHT7hYFFhpj9aWiL+lT8V+2
vew6kRKxroa82R05Df9P8/6Ouqy4vWG+c4OPnAe/IMUTcK0NtiDGsYywqPgqdBPh2Q1Zq+2WgWfH
uzMm7gUH1qsfwfW1I+OwscEWNAwMy71y0r5hmbwIfhqJSgcVSKfm28VekAHUee5q7QyXlijcvPFg
rRrw3omz3QJCp+7uXz0NGGJ9I+9PXmCqM1LxKRJj67F0mf4UUbQvkN20Kk6aA755zQ791NrVuY6B
PGIuhxm7I/g2O0Gg/at2kHKA4Y4JckR4aH7MWD9mmXFzpHTNNRaljqshvtioPxmz/2zaMU/J/NGv
AqAPBCYICTulqUFYzfeITOw5dJO3ft8O9tLg4sD+6qlqsXCMUcsduWiqQ6ARvUOMxf998hA1ifNK
CPXkHlDlJEWbuiy10odCTuINrn3J3zadJ+I0+TfFIYKwC34k6xCNy9NZsxUre++1+7MIZiddplIE
6H1cHET8LQWPjD0OCGmCGi2ObAlJyn5nXd2FAlCTHsKg3tLYUfzH8X5EKZW2wAtl+vLZv8lexdig
Q0ao4Gws5FDEyc4k6dvIsvIGKUhnLFffsjQbu83HqFimf1KPmOPsZ2aiteQAhzKAB3yDDZUZUmUD
7EY31ycwsNeq1JpRdQYoP49hx1I80e0b4ydrb5bEK3zePzCd1EJaNQPn/NjBncoI128VdJ2Vlr6C
ntIR5BqHMYRrkfp7i9v3gEr4TiVr4+AiV8jo/AjLA4qatqnqxGOcNTx7/D/xcrqFTy9v92/G4tkm
shy2OEHwuEg6L7XpU38Hnn/pEk+5EDMrvpLS6+lMUyBt7SJRtnvFe1TYJu5HjgToFej3r+fCGRIP
Y9GrLOyM4s2WXC2k6zOrOMxcmEuMfCnT5kKheucR9JEEdSZ57Tf5Rk+dUxMVlvMPKg/43PYNykpM
rwt+jOzedp7B8muasFCOP3wivE2RMttnqGIVFBIkKM5cI0JLFfkSm94ZuMOodU1wObAZEfrB4Onq
qtPGi+z7xhPfihEtTChbZKkCxhsIqz4hfVzxrEoAUqd4donREbadGSq+8iER+gOeNxBwxrIfz62I
1twxBSijTDSFqWD+dSfTIQvxn9zRKQUe1r37QPy8zLHlagspHCCdUHxGoQLkRpqPyXSXkoXg04Sk
5WMncozKSN11mrydHyJgUWZhWddSwyiVFnonmeTqppz7JDQfD8QDOT2Kdm310hshwL2/X0S0x+DX
x/oSRe4uhFeaTmq2kx/zgUomjNuEEu6VCLWspv6OasFFYdm394lto5ZoTJyR19XxKuktzuaKEiI6
Le71OG4GvIgzVW5u7ys9TsLM4LQhTCvFf8fz8G/z3KnLHUJ1cOl3AZLv5H4o1Y+SwIhXiE3cimUN
KCeHSGeupaaMW3ElYtpW/PNowpNURalbUIzDQlyO9TG5PV+xb9sjFL9MoDSqT1+E4wkJr5zbaE+H
CfTEJ5WgfwOTC8XKeAaWggFaXbQMJhUkftkBgrD6vjgEvUtgr/2bjUYHN6sIuBrp4Mz8/FzLOGtT
CHj204+NjZDidh6Pf0bu6ceCwcs1HA0Ixr+3rHcfKdSCYXtZMGOzPH7yry3mE+DF1tzaJNVNsRoF
fvbuLCkregR55kX/eYU+1k7m4UWLedhhCpDkIHOdqLfjqZHoaNb9R9dpqZwdjLUShlb2P7Iuu+EW
GR+Q55cDjsgWvvHlujLT/N/rBT9ZjlH24q25jLjkprF4nI3Q7Bt0Y2/ISc7EXPo82JMXXn2R8wJ/
aVvFjenI3e6XuiTQvTDUB4+1mJ72YLiDIzwTYzI4pACtuUII0Oftr1dMuuf8/Yxh5GWr0be4RUtf
uwMzYmR137cXZA+TeCJvZ48Tn8V2i7K71SxE0FepUQVYs75QfEtvT4OAU/8n7v9DlrHvLV7VNZx/
d8LgaPwGP83GlpR1L72i6WQ4gLmJ0Ku6TkZYvXcURUtInqzN7+dFFHpj6Jbhy5kWvdO/1v2jbyGR
UBRgO7YX1/f0SJsaJIScfT/yj1CvNXo/yyqBdXFtRfGviECmz9hcAPmQJE8vbbBicSh8RylrVuPi
eDXDCNlbzFpLtl6KCUP3zCyq+h1Iuhe8teLZCn5LnGcRKoNczK2moHNQt3aRz8bcfqcG1zqACxju
jx77iHnOOozpzfT7MKNr7tv3NpTYmixVpyqAXkR5L+MnxcnYh+B4guhgYHYoPhZOFcofWp2CJDjR
k+cjEIpwPZBN3DAzDM6nLbuqJwqNhdVSyD38d5spnwCcvlWliY1Wa8FpuVeXAtJUB85GToYAz/Ar
58tO/qvjd77QvQGjX0xsQnTLk/bBAeGvorHMEArC2+G4k01gyCcXaNtKW9/zpB/sWEWX88EUnxis
cmdRNumOFaibFKzHM/C3s+gIYp41hO8CXKw150ZLErHtmpWHis3bc18nhtxAro3iEFFaaMdehwQM
x7l40P6/4enNeA02tX0+LwZ7T3Q3BciCXHFdiTL0U+5P0brhI9Y0oPrfsFt91HzDdooc0K8onSL+
w4iByoeQo2kXSNcH10G5Rc5ER2X9jTRrx1Xrjkm2zn9PB+6K38SJOoojzxVBocaBgCiBmnfkIs+y
gI1n2repXEA3nBJItkPlj42dKKXv5DfpEChw0xJif/DZohafo+yLPnbtA9SIZPalsqTZ7M6FnNsI
6xKzI4d8iK6G261zKqFCG7wWyFYQ247XmH76Dw5AZ64uwGmn5fNs2j+lSCS70G6arc7Llq/vWbGE
Ekcf+KT4tQJb3fhoeNZ4leeKXOFCO9CwNY62+qWWII8Fbl6fh2T3wSP9SVCEv/65f7rJeDecWvKq
kBml/jCe08GwyzMtHSxQCTMNyM8JAisthuiZk/aWDo6lHRMf7MBe7Skmb9V6tdkcvnfbRK73TiyF
70bxTFQKYzlK5PBTxDdkA+2jsfz5YXKI2DhiRxad7FxxTDsrzMr1FauAgRl2LSVl5+gKCchp3vz9
CQHr22ZZaSKlastJuiNCjevsnWIN/xMsplDfOenQ6noegxi+A7PTQPd6MhSHtImbrnIhxmB1tiJ3
WmUzWjLlmHFKactlYh4LfHE34uiyceNjHsvVAOTaLQp07zGZNolWXAbEvg+xDnLuRXVxx3+d5+Pf
WO5nTfJNRyel9Sno1dI2pp6KrqScENNKfZseMMxLrmym9BuVMpocdyHWQQ0xg4XXejyO7sJXgYBx
NQ4CkZ/J36+hZzxlMQrBHNeuzPUD0uD+yfAj8ZKgaRUcsiRZ1/6cd+l2vRBOB80jto5d6awL/HYE
0SzNs2GnCrI0YGB6FfewYf6XqFcnnvGMTxqgiKPxYa8faFz+a8Ozq8MpR79ljWaex8U5GI0QNtkm
Ao4et3x9uXeQQBtbjwYkc6oWsFDEwAyUsGycHgSxL+QeZmONnYvgPPo+xZOr8Ijusq+b3tnVY8kj
G4FWceNJ/mJ6pdagxlaF/lguIp1jt+y3mLPzfaJYnJElTVGELFTlZZaeNcutLSv75m5vJCUsBRqe
1iQmavD1erTs2nPpNFdMHJJRBUpffqs8B2Sy4I9xs3oTblsIi2r9ZN9997+ikNBn0AjaeOj46Er1
+RxCfydY6iSGYh1QmaquHYJIa6gbWHrA+U8DAeoFx3AmdtUoArxkPzHFQwE8BNFEq+UEVgub2mzB
OdA6PObI4Tmo1bJmvikn36Vlm8vANYBv2+fJjuwv3raqAkdC23Cxl0RzyOdQG9DEMdIpqhGtGs70
1Ka9pNPvdQTvtj8nL8uF2s1Z5UqfJ6iCXj5Ss3qU4gn2cjhRdBKI0xsdp0fI/0WhMnWi/omXneJE
PxuRLAyyvyiZk4TiSAjiok3mjISkxGhGj2bCJHcMEePXH+5/CN/tc2tkRrdMDu2jY9BueEw9etuE
cYuKPHulVx3dGDD2NVEMaLxYUVQ6jF2NwuIMvmOvG3Ba2lZNEbQnwfD17BsfTNxvi7nYJdVLiRnn
2dtaOt45EZXvAURDaEZXJX1ImkZhsVIOhy4oFSn71Q6pyt1OcHKrGAzI0sb86knzQSnC8NTjT5GA
zT5wwGMwM8sq5VGyMcDreoge+js1uYpZyd+YcsZyArIuYR/A9ClTSdMnepOX0yctVb3qQY3IIA02
xDhqsUF5CHfbMg1VWXr4QS6gDkgaKgPDdoA1okovMKchKvIeKtn8BhYpauNrolJmR7Vlr6ybQS1t
SFh6zGVZzvui3gsejWUl6Tox4jXjQQP3kO4uEc4VY23LDT3ZvqDaG/yb01O9sIPgXXB/7p3hW/Bx
gnv6Unhzmunmaf8w/bIzTjDP2QmNYbjy7Y9gIYu2N4XkGqurWJ+fXuHwnQszL2yK9w4+VTWR9gsP
fEHYFH/MoLY1xQwBg1fiZED4HUnno4wR4dyCmxaMsw0oUrKEAqXydTorvyo/uAV5m2uG3n8nlzXl
rWE8Hio1zdbtiz+hKAFVp0wQF0dTTUpPRWGNham//2yxUupZ5i2F6W5yajr5kEG326jOs4mJsTBc
lP2KKLNwM3/Muv9IjyVhZEL0lGmFl6LLmZyaB+2D2c9o7ZIHOdyv14OiAZiG9qb8IHAOTMXzmp3X
X/6PZS4UiFQmaGH24oklqpSvgFICfHIpTQA3uudUfGCLjl/x2/SZALgH5MBduyohvSwHc3HWnIlN
GXQhUPUE0Gzsr/R1EmwODURJGD5Tn5vImNR+d1DJtFYfV8XkAcO1dVK+tJkYPS8R2Umv2zaFyHFW
LD4IwQRzg7d9TBfc3IasCj8A9ZfHmkjlmQW2Wh/NDSgbM6sGloCH5npWAbg23dHJAsqdkUmSKk5c
/is38nH3pUn6bcjBL+hPH8pI9565gXqU3w7DyXIiU7buI/kuz64YXYKeaekqDzBkrwa2HZkvUL9a
7AGVBRbenq72WRX6n6qXTi+ZPIrzaSzumrCEQL+ovBocos4cobjrCwkaw1obX17dt/WktnP/Y3tF
i1ks1/d/mBPF6oNmDfhwqg52E+jL157jktfPLwDeV1tzqeVRzJvMtlhTVlglLGbNpdSYPyBe6G0V
8bk4PsU8jyszuM35JZpJXXhEllakOraodCDH7+AtFlu7L/mMj8ORmvKYEgwMm9zHlRDGtPhutE8z
0GSXVdPGSMUBHvsUOcCmAkSx4UhyWiMZvtW6g+b+Lt+mdNVfwHNbHPm/udTEc0Kt+geAJ6s0J1gh
4JdgzHQe2B0vB6e5/VXXdnI7yP1pnysWAZ2EkJHmKL5v0BOGn26zql9qO0ccSMsW7UWCNj6p1A3k
l2xQpOefT9QxZnzsfjviV6wWhY4pY47nmaD2u6DwBixoTgspuq7GnBQAUXQ5apIkHPezzxZWceGD
Ze7xT3z/neMFLSikI+F0pO/9Ev2zjcW/282/KmcZzHZK6jdSCjh7KK1TAo1/zTNTh59boG1GdT1c
J9y8jCNYUuzpqTXZyvBKJqTCtFpC0j3UkpzlEEWvWhOOvE9UQq/KByVR//YDGAlJB8r1rpElJOqf
nLbCEMQdKUO2I39+2QXQ2MWqEsrFdYqjnQauwoUlQjDjJCe656OldQ5h5z+P5WkwyoJa1SCzwSoN
posN2k7lndmMzktHbTnbMkemK6iibd3na3XB+V7bXLPr7aBlYB+ZRQvIiWn5/jg/6KWHgRRAO/jF
Yxxxtp+pIH0rNChOw7NZeLmYN4LJhSoCDkXjv5sV/3tJusJ7vJxJ4xVlmHzHwZ5H5NRQVXCZw0Wf
QvhRT0pYyxlNBK9Rsj1VfSPRB5dlrwpwzMxE+n2Lbl+Oniu2U6uV0+dpNstCWNvQVGyYBdTNR0a4
bNpjFJ7HoupZfcBF6xa/8ysof+XgR9+XkL5NZ1fmkYcWL0rXTuXcnfv+pY2NDExk0CIlrLCWNYcZ
HSCv0ThgwTqyTi5J/y/JES6kqvYqtdBWz4H6ZWk9c6RieGz8VZzDCy/VbvVfKZjg8DtH4Z0mYtLz
NYgBw5FEUngbHMTwJW1xWVQ6PkRgFl2s8pEBVsx3tOL6fy2W5qGDBwp/o3dDj6QZEMotnXpp7V4j
wUblHKOGiY1WDHNP2mcSBO/rmHKonJCDYEFZnc7VKJh2jHCi79MXjCf96oLomfXULf7nRwjsXKS1
nqs3GWBWgKiq1qR5AhHzrNRecj0oALedTToNFmM9hbX9krTGnav7G4thD2WeBU58p9v8eW/4Lsgj
NwrLvTjoi4IORDAhhSP4Z5RkURbbh1x7KvxSP8SKYjBJmSVnME8vW6/yENBQF76aP12FsULqMo5G
kffnu6smLsQIPPErPCsF5mO5BYpnO0Asgxu1wj0EarGrS8vUCu0Qfe3e78EnMcsUjYD19W0lk34m
wYrjAHnZM8f/oz3Ni314fLgoYYAkSz4fU/pEPXPW1OHuoZBUTh9FiQS3xISRNI6F3FcrvnouhjvU
4d6fMQsbN4Yp7xIiIRhsd69LatA7jSjvJxl2Ut5cn6oG/Ob62Ie6ugJo7qMF/RGjnkq/6Afzt14B
pN8Lvh4Kd9kE77Fepi9CRI5yQ+2wWLj7l+HpUsSDhcpeODxYT7WKzvcMLZlA16vuZtVIgl6VpyxA
EweTCnGB3b/Eb+5Z4il/4Tzqa4BZMLJMqlp5UdB92otgZllz7pavbp+CXXCU4ba8wks1EceyYiTK
qC6WWP8lAHfAc71VsQu4FlAixccGlmcVleH1iKhWPOWxK8Y23LisWShhzJVKmGIwf6Vkkq2tixl4
pblVrvX6KZYIkfDcijOcR5fM//Uc6eQgb57P/H9QNmu7sb2hFmfuCndYOXLdr3mfZvoeiDF0DcDO
QKi93Th2hs6IVT3Cc651ZLVzblUlT7Gl6MmqSPKzgbVYpwOjFtlx7hQXz1c2bxhVqZLtR5no0l7M
Wf4agnFG/pDOa6of/f6PDlzSVgRABrzzeeYgCYXgzbUaMkhwfE7X2LA8aRJiKxlVk0Oo29Lkuy7I
V07jjEbkLbD5N2CboAt74dgx3aZnm9VEFBjioqDeG7c0EfQJPK1yBGv03Blfm0hjPjlcnE4KFHZE
HPnKranklRKpLn5P8s66moRBMjif5HtTWRE/qUoJXorq3Ce+DONheUCNIm9Di2Fu6AVoTq0cPxbT
zOTXFerSJ8hLJcUQ5nKFrlclVx7JlasLHJ5eYY5xJ49I8AgNZORmqlDBLN/leBPqgfftJrINs5W8
Y1XDZF0df0a9JtUjerFMjRS1vg7E35a+2UW6jep5KGQD3Q8a1rOEk0OR/YWQ9J8oFOow6BiMDobY
N0DzPQnUZtLGMgvqpxJGTV9oaGuds0hN0V8oDc8j3CR8r8y3U9i41Q7YHce8/4Oy7IZyTMv8L1sa
Q/Na36Tbrl3gU69kuzHtZa/BBoxLdZJiGbV/RcAveZTnkVo6xXTSxvzmmgX0HJTwzWi/CJz2tcmQ
cmzQ5Ao5wW0YBUihwWtV6FsMKFppRLjHrRE4g2KfHdwsWWllLgsusEW9F1fHqwTMeX4WA1njM7Vp
2Py7dNn4r4PGvEk7zv1+zo/I2Yin8OlXqtOrYTVeMJC6huTusVsd8+ZIV4RBEdr94yBEypHtBTFC
S2fOhXW2duo+dJh6zw8+2eav7HvHGNoS/eP5TRzLkAyMc9Qe90Ce5FgMm3fRqZTx4z4rWLMbWDm2
oZE7db0tU6DCPW7XW7Sd9866HALm8U2G+Fu9C4cRZ7mwVwWqKiU7MvxKhXp43kVeEviUKqN4nOHg
KBxION7eOxeCDx/iEZqKWzNPzFm6eVuDwxPIrzf/Fx/Dd+LVRvwBO8IfQgy2uwJw47NaWAmz7b9g
9RSvr+KokoFKtA6jrBIKkmOmdo5GYddkF28uD9qscLCSniZ94tXuyLPia4V4P9D4sh2ZblTVQmwX
Yla1dB3+88lyZWDIP+CivtEVFCNAK3lB6UvSc7PI8nkqK8Ao+wO1JiXVpU3s9VYC97n1XObcx8Nw
A8+q+q+f4bFbkcU38PleIi6oNPWyYSlyKgJ6/Y8rpdsYrFzwvTFmGoPR/PtgmUugCLpQZLdYlGb5
UO430OzNg5pTztHF1rSOLFjbEkIqvV3eI3wgCN0bBxjjG3y7R+wn2dbGCWp3dixQ8K2ZNXhE1VyI
P8bxlizFiTp2jbPSAY9nImJmX/Lb2nf1gPbOga5uoiZ0n52k21H2fKVEX2sNfbOkcLZHqkeyxHYs
umE/kfsSdFbA8GBMm/zWiHyqecMQTqYEjan9I3nLPIHHHHChPbaFBhltRgzmGOdzmwJu4FvKUoGS
nVThA2Z4NJ1zRXHIkjABbqhUIgSxHrshB3iBUV3IhPSHsTxBAtKnmfCTCCsuY8COUdm0Le6agySz
zpco0Au47c3TjfoJSiwWCQOdmkSWxXfo4m9gGf96RnY/9mjXWHzIbVu0rn/kJFDOurl+uTOM9Mw4
DxTQ+y4c/t4tr7r35lslmBgXKoMYXRqqM4AnA4HFHKuVBWJ0jJiYVUsirkzILlRm8wvvH8j4uzUA
5/eHUXGt3e9TIKF4HT/xnvXK3wQfOW2p9wZ+UEhHl0LNX8vBRvN1C1jlCe/ciTX9ABdRaC3H0SwO
EbJnT3HNW2mRhWYnRIDteRyOta89fWjYO7HZ5jecRVmC5KTRPTedoBMgjWQokhhZad5fdvU8OJjJ
4UbksyGA+HSzmqdOSAzQ89xEPBTaHDUDi53A7IQYtRBj1Q3lzix0Set8w7gw+dOWVxAGaNEh9M4G
FbIjZQxZiWLCJVHDVrJbfHK/TOn79H1wvmmEjsrb3/OT39r0pGgSt+Vk/rkDMgqBTYTX2wA6SHYp
MbAw6Hm7AnlayFjmm+cSw251jy1fPmNLj9gCVgUBT5mrbR2tflw06i63A1Uc0reTZxxU0eQk9G6g
7IwDbMkTUsIHOFQhsyPdlKxXNsPfcTTxQeN1Uxtd/O/fGNsMowud4ddQImAAYdUHIcfaY2/QWe/H
kR71aBoh+5mScqUA7clPF+PAwnoeNGpSi9I06G49h+5EFfJ9zV70M6HAhqh5TbtEjDKv23/CNBYe
iC3Tu3FtDFFpIuuitcDZIeQrMqLxWuoBVoTazbtsfTDrTfpX2S9o46gsvNde11AFY4t/dtnR+sWa
Mh3FgghGQO54f5VHBaReWUe1XAdcSAKjwOwMEEl2gV4I71HFO4ywEajpvYyk4cHe2DlsjKyylnT0
XKdgydFIiluNaNh2h12k6ErTz8zwP+Mtb9ZuUg0XxHQjRNmyEMUhc68033yUiFP4+/CRiJHOsHwO
ZBZVpQorG1LPI7XqYnzuu28Q33HVyCKH80NOYTGH0nq8ayVXZwnMpv7mNfNPY5xF+lrrZXm+Kg+B
xXHy/1STWztLr6R9/lmvu833HqtD2tC9W3LHf/YISdEyBP5oOk4BqJHEYhqdP3KOBjNzTQuQZ+Jk
ZPm5NWEOALDP6sQR7qe7bjLi+Ba/5YXdV09F0nU6esK3y1H3VR9mZuSYfWSAupXGBgCuNsrIU/qR
HrljSb6Ub3MLrXpIyjKunLprmlLVgucZCgxv/bBfDMrJQDFn7QaTULUrZlWxSSP+o8Sclp+VkHZR
9QrEo+cLHcWDwDVn5PheSJ1zVH8s6VFQ6ryy9zlhxNtSMDGU+a50W+faBDYxhrXGudP+amEcMrbw
Ov3DJbwguhFfPIrl2utFTUMZVvbhJf9oZpbA8KVE6fTfjxX0dTwxKj0Bdia0x7FK/3jGRQrSQJtn
8+sWAlaM1zqs5h3GTiTAiTn+B8Kc1q/zcoebPAj+yis5yjalUthyP9PYWVRun/huAuX/bcP6S8ZG
D10wZyRFyzJFYD5ZwDabFGEgmt5T0YRcsZwkCWg+JZWEBVKQi4q7P7GtfbAI0dvctyOvZ3NTICxX
y5qZNWZjgXZpQnoc5NnRqrhh2RlSdEsQk5vPh1lQ1F+syJhOhd4d/3Flgk/8768BvCNYjZ9r94K/
R7VDDoIk5mwe9x9BN5fUR6MHxcCZ5bgM3aT2pVzSVVuBEM2U/2ZeugBA69RgU8qsARSKzZNSKRNs
D4nHQvuV+ysdPBYOsKsnvh9nnDLQI20LSOqRE6Sibv89QBBgvarZY5jZVxAi1Nv2ZEEXEIaeK2bb
LukrA9CO5oTwqGO+1Ci0RGc7zhtESd63II+AZyXvF5Vuck8VOLFOpj/4h0HhVrUoFN7NOL/YzW0f
2WWk83H+CsXa2bL9Oe9IqXt6gI/vy/1sDEIIPrVw6E6VmWOPcuubb2iS+3GSMyaSC6FF6YqVmQPB
MFRBR38jGWrcC1QfrCgGxiOfilccc+WfraTTrqiYCn+GDDhhKe9xA5SOF5J5cUzHWCqUFlpoOnf9
Wx9+9rv7w24x0If+X1N4/Y2QJTzFD9ND56m6qJmQa1jf5pNeF34ba6OHaadaAidHcBiEn0xaU9AV
SJBm4uLZhf/aZuRyJT/z87JhdpuENFro1+xDFaNDGiPwIvEnfnXE9wxq66rYNnodIvzKWBOsrrLO
+L1j34NmAWE0OR7Bt7Gk29HB/rHXJDLTPNUc9WpRgXPz+IjosGuQUIDjaadRS+W2suPRdskoIOxE
xTy9IjYf3RmQvkeM9+7Wsg+I3o3r4e6D+1Q/ZtP7emQkgGbWsPCkp9XePswjBX91IDyY2w6MX6RZ
q0fWtoJ2qZ11ULK0L7AX+taZpnBCdePWIZSexycqx6h7Jz5VxQEK2/EjvN3pd30UOhYQugyiqql4
vvgC22WZuabrdM2YdsjgiRAD0brAeEIoiGHtj6rtd+r8TcN7cHtFpr4gbSrojavGaHx26QMWuVHU
M5zPX3wG7ZtHL0iJTwJpVAb37wGxYUxK7/o9YwQiiL8Rhq5NaKiJaFMwEFn7vygN/4v7u52C8Jr9
w35xDYO/6f2S/z6OouRefPIPhFNSH6Px62xci17ngRIJHx1QQdZZtyjb7u6Lpl1aZ73lbRgABQAU
YhUw3IKZbiD+IlcszSIuOKYbEtR3zQP8EVq5aF83Cs5PhOJrgCkE2ef0eaR1CDL7q6k4FlxAZTgP
d4K3DVZs0g2Y9bGClVY/PasG6AQw6evvbdVVpFzhxusf3gUS/32U2afGkNTnvPAa7S1zQGQD0O5f
puuezWcftfawhhibonfsUUtUbnaSYO7jICNLkCECzTrqrX1Ojf6p/4/Vk45FS5Ae6LHewAKH4oOl
bKaXiWlCTv/rtMEo2ZVpOUB4xI2kXObECdMnW6+ktT6Lv1K3OPmN9+kYtU7TpAA2dX7k/MTowP0h
cwgdFllghsM/UJMbuOe34J7hZBIibNJ8tUXrtQmQ6sMvsNevymAPsycSliiUh71UIZrxT1gXbTqg
SjXwlIuxyykLC10w+ChIYKdQekIApsespsEQow7+8Mpsk6voAVHV999uTpVi33R2hXN4NjROo6rP
hr1k3AsF/bT3JQa1hzQrtkFLjQnpUTBJ0RrdcvZSpAlBWlHc8lCjFYXO2pLDqR8UfeHnsPoAbDtN
AKEZ1encpdHocttlCX1tTuUhN8WUyECmGdCw4KiJB3lVPQ/9F68BmnN9g55gQO/eUerLi3O3eLZH
vydgjCUxtyiKA23r0dq4WB0sYtfKSJdezq8xQhBHxka91pjZWTNCh+4PFJ9qf7BvWEFRPvVO1Lks
cPrD28L+wk0f65d2obYKo0538D3v9Did65jhogAaJQN+5QdT4hO+STMA0l+BT3FA9SDFDcBtl7Vc
PZGrOdO9538ObY/3ipnTSfTYPkrxhqAfgmlO5uBa+y0wQybda3swomw+ENhLdMRlymhXivBUaHxR
dOIdm/ejA2nGG8N0jpS2zN7OiO2Q4mfesoySVEiOpd9eCKrBOL73DCb9FPOcjVplI5ZBVdI9UKYt
a8lwUAs0nCvO52Sj56a9bLvfgmRBEIdkEbWsLLSqJXb67dR2wyHXCqur2CeDrOVdrtk76YUmkdvM
qUYKU0u4RHVf7O12yKLUrrHzVxIxrDlJHgwl/FC0IymlbelOO8j3KLyVHhFTqXnA63vMmHorrqay
yWXHaXetjtyhkAwWscQln1cfIEy7Hmjun/SxCSWBiuYN5OMKlBvrAe+kzciS2fp3ghkkQJ++fzBe
rpf9KNx0DZk1NVO+0X4DKc88ooUSI9/PAgao1K0L7VHqudn4MVHseoaEe6xnj3L5ML0FukUf50uX
uGcplIluthfvr0KNxnEaFkNDNH6S3J3ovUqsm9hj+Io08KGQNADTI+EslML/6tlo6dcGPQHGoWAt
ccmUuPzsJUKcgkCRr4q3I6eHlQlIWXyNmWUsBoJcBrJPADe2WynPVN2UnX4lIJTpRaTrRsZgH+iQ
DaAKliR7WUlV5Ry6KoazmYm57WMNaXsZWr4rtN5EjdkLW6vEySDcyqqwXNbQVuJgJYT24QBqnDVi
nO3qYNfqtnTJU6Y4qdWhb8nRZuwaaTrlEpD+pCX1KMZJp4ukaBc7GnA48iFH9stPkBFt924Ul1yV
r8Fdy59rkR3shXyvikCw0nFwht2iMpZtH0eJOipuHc5SbxBHNRubOY35Vd2CwZ/Wi3j4ujVnQsUC
i3lj/Z/pcU0ORaZCHf8zwlV+FVOiAjCk0blIL4D8czugFNEsx4QY9mfpkgKYLkkBmfqjaAQVU/1B
M3YtRZI9ONRvwQJ8LyC8OtGNjsVi+tg/GjvYiyY7Tpa8uQF1clcruytPuLdkh3ZeDvz49YZtngkb
iy+EQrQplHc5aa2CgHgzcMl140KA5UxSWTgWe7dpKbm44ZriRmygwWX3LFOU00JDQvdiVUj/hlGW
/NKGHyH3LOTmudHZz+33oOKPGIrgTBJap0RCiGODrE38U6Jzj6MA0gvFDco1xJ53eYEVuPBLy/8a
hnZ9GfqMjjrXEGTU4soJQxX7TE2cxgBQo0fhNydzMsJoBiFpzNsUrCYKamOfJfxEqLE7jkBrRxjS
cmvBkZ7GaLY6eyqYT2DdzmUeDNa+WhWCvG4Cst7GZBLFvmVe9Y4eUrr1AxHtWA661W7asl+3eUMo
4DvGBHole01xciEUsptTW/K42vHfYatLnpdX9aafcS9XGDcpFgyaP7Kfr4efsxSIq2dPELlL5UKi
f8XhDYUCuIdUCCPTtGIq4sbUcYxfJGa65wJpi+iVSLd7f1z6PJ3UFYrwT6tATm+1av8LZrZW44Er
r6SBNB0MvMne7OaIOhuCWjQWa6b5YJkBC0KmX1qIF8b/D5KXMopSsqei/rcuIF2QSXeY+czQa7YY
MqNXq7kaDoRwOCUxGLLfC6W3uC2vwFDUpsOvP6aK0AujpBRl/L5QDh2AAOrbX0F5GAJW9OJ3oAgF
fek/L/sLt1gAOvhK+tYVWO3sNbykSLJwTEIOZmq9SyOausPORwHrbVuP7cTIqmROOTDRX7nQ2khx
g+Qe5U3Zru2AD5kmcLP/2ZbT+IIv6Ko3iGnc65gpHjRV8yTVspXm7sQjgnAJO8M7FrwqtyT3NW3a
iRtMdW+EvKFpWWWAE9hV8HzrySYKO0k4IQ3TMz0+MloWrEV3qMw4olmc+FplKE2xPxOZ07H9dNfj
nIW2hsmLM+SzjPNgiBYYGBnFsfzX/wR8vdj3RC8eXyZpXYDZHRb/rEIg+5Yy3X5J7twGLsqC4Y3t
cjQUXPtb344PFSuw6sw+8HtUvbsdZG/mPvbHMBtpincKYxdZ+yliyG2GG9TgROWoYlpLJKGSuNdF
1wBDAls6D4C0bnvqBxYc5aLNdCFwa+yDKpO+eMCKhsaQWGFDgwfH3xseva5xOb7bSUKxhEo17AUf
zmIZbcGwivUTJhKoCrVOdsQwWlsuph3aQDKF8V40ebFYb0N1hfiwn/6AtxbQa0BrdCmbPjN/cxcD
dCANUuyR2z9vxvVFyY8jyZ9HkLKbPQv5xb/2ru4eG3/F2NZaC71AJVo/kk7sH5+9rT+EbytHN+Uq
bpaSCR6agjSpYBLQXBGHQ0q2cvT7qm6+qucLEkK9hKu2ihOnwTIb+AtyfEuTZCbCdxO9P/ti/Dhj
ShAXM9u8FnVUXqJPRbcXE8QGHiS9HNZiGkIM5aYcpaA6mThJHyTo2X5U6sxlJ1Ixoq36n5P4RrnM
bvSvP2W/cwpFWfA+mtK1LvVjlWP3tcnIDDzJv2g7sy+pRp1fpPq6TWTI27TZWkCR8Ar/5ZLjGiAS
1GAQgB48XE6xv+gm/tg+/PuNbtWdS9fU9RvdD3fgbtfnLfHqBIcML702NuVbeCv0eoPpd7snbweT
PqKCta+IjD4NnaXmosUxSh4PjDULdTQvStn1mCBIhCxz+6XDHwtKjyI03S11WfMwBIRpZu7PxxBV
OWNKIq0VI+KlkHK5Yeql6ay6KhH1n2K7WRI+9l8pmG8PadtB9brrMoULWskLENdOeg8g4wLvX81U
URfmPW7+nbQ+eQsUDhQQg2eGfai2TmzcqYi9Fvx3+pLni6q8fTvc5U818TdHpd5XIR4iz7FTnfc5
PVoqBgbYoCuEoozcqtBNceClz+saKH9/IP2C3eRuwYmIc9ErV7bFiVjRQSx3Dp2LpWdgU13WDB1b
qr/0x5KRjkqifZw+4QLbo4OPCkmVm1gom2QFOD9aOU0VVsz82yl02joNuqLkaZp3xWLDTwpS/PHA
nhAgO3l2ODlTcb9W3zSLyk8vcQVOKs8acr8ZvEWjkBEmRuprjAM0Z5AP1LjPdgT7s/gS+QFW4QqJ
CROP8VDlcBRklOOn00yI9VsAzTJGz7ygNzeNzwi9l7RrQPUpBhWgP9tuiLJRvXCq8jaKqR84VCnw
qG4dD1DfN7ATd2yfP21afKy6/P5t4CUxVA4GIMJFcQkUJqNDUMKT/whBBWtpHlNvCPJUCkPygymv
SIKUGioUWJ3JYIGeMbhLqkUKiWKzA1XZDOvU/H+kT9ShACrxv2HSlQfuKBQF5OkrAQnLkG7/IOtG
wxoHq57nEFc2/xNNyyd9m2BpWFkGEf9KA1zjedxY1cDTJ11R+RqFM1kL5wucueauMU3bL4AEON6E
qHr7MPEzvU8WWtNOgbSzL4TreyYroCVY7hOOB0iE8VT8pbWjo+6TVn/SYIK543fDy3j5cHzLqad/
cxoYNUvxwmUmi3tk0YmR0kFZDbKObO7bd3EuL3XcDMg54oiifonjPa3l53QC5Q4q6HP8LhqsCOO/
9DvlLZo+a+ttKnvcVBDAWFazbTjH+f3DDxIt5tkVqp+bWf8ZDz23q6YTV96m3AMTXD8/eWYR5mL1
Mio4sZ7WM/BWjqiuEDNKa3xqdLOOtX/AIMwkQayZL+IuePEm5wHvUfjppZ0ODmPURNSEoCLx7bRx
cLe/GzUtZ7/cSMhDCMJQ4URWHGspFdbKIfszjHAq8wvHbl3Z9ScJ4wWUO6PExlEVkFDZp/lYVEyv
kMs6H7XwVXWAYNkbhWvTjKvcHAgLoTL2ucXF3JpI+z+AYf2Tq3KpoyTAseUeu5SIWGwdY3KYZ+Ri
vQ868NuezzqU2wyQGWB7+27XResjPKxW6IFQEpaAXwSG+uNfsIB3PMtEAWXoAVpv5mJoOeijfmly
BmW6mKdWR1IlpsYz4CmTo24Q8y7LjoknyHKyGUSk/WJTF8SJjgVwIjw57ADCNvTGR9YR7Zq6l8wK
RfMpjKBQ+3zSyWXmzAe9k7yslILruGM/aRU4mHhrM51XrnyfG7yk0YUSub9iIm+lwYCdicr414Tu
Tpm1gw/2MkKCiO8aXgIE3jEh0hb5QaDddpA2UHryMbwGpEe8N0pbxNnDpYvtDEZsXq7FzOh/zMJs
eKsIkEw/V/57dvqq+zPn4pUPrLYo5vO4xxCdPvnc8egwBrLPUP7PEA++vVy1AJme7OY0G+qcpQpY
/rxbv3HkXrICgBMHV3YbwIz2e4puB2BaXsuavlq87obHIpAv1TKTUxgJ3SAEQiTE6i7wxm5Mf2P5
fxKhkVWumJqbwuPikSVWtwh0s/7jkpRGjwzqCPsHUDcMWppT9OoB/OrZy/Yi9vztUfhe8wBPs1Rw
8V2AL2vkGw4OAMVl7Cmf2d2pHro9Bh2+wo+asnOrsE/bPNpzjMRlCzbevOurz++LIcH6J9AwIvS0
L3UXzqnQ/enal7rjFptgEA47KwRwe7DOUClYzhc2TcHvKShtXRQGx7Ye81A11sJYSRUyKxFU+5ZX
ohAaDyV5HqLZPgK2twrzL+2bZDhVFLT74iUTPD9MZbvT5Bnwh1OWO3eK2wKgr5CL35+3wHCsl+VX
DflZtBQTETN2IVkUOJOXUENoTyNdjrbpzbYon3BjxCX47L1BxEQUIwSxwtMsuizLh933QHB4y+uc
saTpO0Xa50Y/2Ufo/53IAQeUH0ITKHM/XOQmPmc43A5LYZeh/kcYuooBgzv9DbeFl3a2mIgIcROn
FXX9tnDwwE8JmMIkETe9FiPSELZftsyi1NQm/g+lrwTL2E6JVcBkKNiJZx96mdkAvvaMnsaJWM6k
ABdVKz/idTdfMTrBTz+0ptIuOjmxXI168NAW40zkXXYjOlVMFlQygXGPDHBR+iy731mkXiJJlAHV
grhJOox3Lcrj0dtdCcAwMcrmyNaKv1fD63uF1UmrPdaGDudTdNM7JsMcevIOydAcYhfE3Bm2Mk9V
kIlWxLweCYq+CVffeAxPhsS1AU9fr3Ok4OXZiuJ1V4pKqVtGP8iNyOvF4vAB9TW6QDmA9Ot+GE2S
Hq3zFx3VRpxBzhXjqOSBY9sbqiGVdzXdAP9qG/XlT6e+/OhMNSLQ6VzMUSTv1Wl94hB4fa1PnmUn
16HzGDz5mB457GCEx7cTyrBWOqvdAwVT+1WbsZofj6i04eDcE0soLl04h6/56IyELpa5oqUIYuTX
Wf7D0fsa+qZCazPqRlqRLkEGScjSkv1dVGxa/iZZOTHCC2NaYn+0AjrkbGL5Bes2wU9eoR1w2uLe
AzWjNZ/Ji2wTvlXnXdeZ7uUcGKkHnlE2Esfw0Ezjsg5lnI+g8wNlFLiXtarTjVkGiZEJi1po66ck
ynPs2F9a16ns4QTox2a7orlclOMWhF+jlMOScAQeWQRWUfjGf4/aAjpmHL9TdRbyjhXkZYUqglLY
8z5EkM1RFRzBHspC7f+73q4gb8RIYIuPy516S7M7cFkk+HMB0iIBSWxw3l20y7lD9niFilSAL7LK
Omf3gyX+9rUCZmeUDhqej66hvGqgpQ00hiS5mggAqQuzFVgRCGkN1JO0YB+pXbor2rVbU9QJusbg
3vfZnsboXhLPR+6aVY/D5S+JRmUhozhw9unPOTuh4A8i1/72SgesDUcQ9paW/khYVrS1cYGinBtL
v+PMfl1hoL+e1mNqHn0OdzDIqOSI8oPTdsKyQ+9ECD4w14Uc8vJyyGz48rIMyYbQhJeEyoG0KYZO
gSH8LSs1448iMVFsv6G8JgMT/YfUAkpjHherv70EnbZ53vVLCiFxQyvuinVUWV7YnAyCQ6TjXrS3
ElQU3EzXC6yI8IZbvnN7HhxxZ/VLlBVLCXC1wV5dnbUfuih4cVF7gOdeyj2Pmx5azJEpht3vPXFo
DdSfYzcfyn1iJkyrG3fraMq77NHGHUolzvBgZUM5czU3tpGvybsXGfjyhaXDx34vVtEzqiOPMV8I
0aMFHyryv8nUJz/QER2xeDIY0NgWBimAtJ+q6pg/qH+z3zt6ABg8HEtPjDx9kniu7ICjwxjkFzzr
kwkcuZgF36QcM5FjaROBp54beiOXmHfy9b+Ffqnro1ApjW+VSXIIRIEbPdyujMxJOWXUM72summb
gg0Gv8RmVdRJgdSEP8daaSqkbBMzNmoVjbHwragdoDck6HgAU26JxK6fp++u9tapQN37WBn7vPbi
TIVgwB4kXY7cBgcXIW0XWa/eHQzfpbA4erfOqqgKjLPXhrK0tGel4oXlVLNqkNBmhHsttKnB0tvP
j4bG4rsXPLxAJ4mbYeM7eiI8JNcWBQpvB5gpM91u/DCqjdpBNWqJD7CLgc9RfO19ZzgU9XD4fYs/
S9WtesBnz+wuJPUMd5QpQw+QU5oaciKGU11+ShRSPYlhw46tvcsObyG/qYkxjJHWqtKZU3R8kGio
cM0E3TAzMB6HKAt0/49n1a6zL2EZO4xtsbZ2XiksF1OBeZugt/jrZ9Urh0zKYffZqrEs+vxafayP
TJDIUv4hmDfcX4d28MwHI37YsfO/yLNME9/nTwQ6V9GSji/Gyvpfujh6TlZt/rXVW9UEDWLvwEpG
DdG9iV5HPC9Y89lZ08Df5ENHooUKeTHwNZJQWwe1I9+7ztxWT1M0QXvu1ceR27nFRbr/yPM3lZCe
GsI8YG2nKJtk0fh4YAgNtS6oKI2sH55n/ATefoNaFz7VQnlE+m3AvaodMoKIb1rR+lZMrUOo8jSW
Gy91Ut+mn1JC/MZGvKUnTOXpZJtEwAnkL5S1OvJBe6sCjBXT1F95TWhrYBPukDd45EkohG7BHrvR
clc45NXyVWFbE/YQwHLZ161c5t8wMzB1jx2GA6NVc4PweIbmDRWg1DD81JtJnBVTo2G/PbMoCN1f
9JzeFrXlZjSAznkDexHV2/VNrx6KpFrlT41C0VqoZAQbEmswPo3eIZeRqIqdwdy49XCTFA9nawbS
S0zAPnOhfqVbhrlMJaZzQQlXS3ZbD+Ik0s4BwNKSrkfhaGCCTQDUh0rCtmHn3/J/B+2yWjoxgtZN
OVpkrVduQy8gfhZeM0mvYcKmMqEccsz77SzTuRxkeq0jyND1bI6HYMBSDW5WP0dPBxM2KHGv9TH/
Vr3Qb3b7h/V81RzJUcVTB+JjpMllKEqppj1DxUWbwH87i7Ojz3Hv64kH0sQ3htHDKeIGvtcdreiO
FiWmUWNmSSPHXQvBLvOrOB7AZ+S1AFkTcbrxKEkdLgkj6ivx0tIv2IViomR1a+bY+qPOMtaFA9Uz
4O+ZIxNefJ0/BzP7Uk6WJjri2quA5nVEuSPu0kgKGl60dcFiyJBPZ20S2g1FKZk0oRRgEN4P/N3m
H0OlpHu5kRL5PFAWFWYxNkUlkVU5tnM5G9xpz7DwA+sNvEgZAFlEz/Y3UkNxLBPaHCvPcP9wVPX2
0UI2QLt8AAfdOlDwBtaiItpNp+NE1fXPEgMkIKCXsj/guRTUhry66GIsCCYJa25G9b1uNVFpJHKG
Pu9nLNAOIhhLUKLOQvnlxS/bulInjPUnTnoFR0jFZ3GcphbSENpjXAAEKYzl+A78sH12EkXlEea9
5GcFQlqVTPf8pfn73lzR7Kh4cghf9Z4Ga+cEyFHprJ3MBGRMIbffDwWMcgap+Bejt5QbgnnCUgCG
XHDTr0MMRSMUvSb3XAXvRUsBykGcv5Bb3vskmj5VAgcbiT15Kuv/xl5SFWyNfv9B/WzntnCjIPB1
MpYHYKpre9+rF7n6+dd/WcbvpGosey7pJlkkeWWpd92SAzAAoPhyfNcGCQFcEVUfhlv+LmqPscFq
729XICeXVMbnUwdW7teaq58phtivciakXMTAGbKTvZCnXH+DYUwcJ9J5943y8QaBSy7WbeZXe6Dw
ZpnyJJYqAodj0c7y7k9j6xUI39k0wPlSflbZX9wSl+i+TAkCt0KJzAMsn8BDI2WFqZU5P/iDsyVc
LsSuN7Lztw1GwdDDcxmGSMds38ri3Guxu+UkBXoKSoSTIXLeInXJCwU+iEIAwt3oQ+GUFViQBYLA
iwpQjeUyH6NCQCbjVIOFfhDOqErX2y3a/8fB8y+TxoJmDpDG0jz0Vn85fBbUud7zaCRqZ17V0/68
9yxZQkdqZnsciw1CdTWOU9hZdrtwksFS3q6OWsCJr2MAO+U9B+zYV8PNNuowePU9yUsuD10iDNDp
1CnipH1DRMSf8lBMwUUP0oOZqee/KAsUqaI9pVYngD3w3tFhCEoqqgOemdxpQluuV9IwxvUG5QsB
DCb3f6Ylfj8I6Rv0aQddAVut+HpluCo9F/TujO4CPHE3YDLbjA9q0IFpPeIVaHuSjcaQH9gGGibR
nnErle3iGmntYXM2vCvR5Z5YOsz/KESO6ksTa1Xh2dxozf2Il8jaenrRWqMkUlqqymaWlFR9dMNM
6ma3cmUAQnd27Z6Hyn7Nd/BGsdK1YJQRjrIJKabJ4p824nw51W3V7q8n8PkX5u6FChTYXlTpfU4S
o6e8/11g9zU+4fRtlmLNnMqmFRrr3+jDdMUT8jTtnr4oo1jF97iKNfnAkWYVbD4+2a+oEuWys3Hf
7dHwadJnpTLOkHh47TZ8dZrAqHGFJ6U5AmdZPAHTj9Efx9bQS/e3H7lUDdGzGyzkclrhf7QFxUkG
vgHtEiigsIW1QkC0D9pHQ5ni4faPmkY3OVTP1p/Dg6fa3fXt7ZsE4AL+zPaDgVn68B8xkp84oniD
/z4Hybn6gyE5+roupYfn80rUKPRzp/x//nQ9BsErJmKxHDqbHBR2RIPKpQq8NGUlRl7q6iCKfedk
XXX758Z9rwUIiPwDTdOuzoN3PLr5hMqBZKLt3Pmlydow/PAbQFfzS6DWShuMxRiaYKrK3D2XvDIo
StfVN6rtxpka6BTKLgIkVI6Qd93jJgwwGEb5/PGdAKxGGTO0KJj/RBWKgABH6d+F1FKH8CdLkX25
eDjx0gr4YwUG7/QuD/lFNS8ujKPTiJRYDOzMiazk+2HEx6j2kiWSCJav49lbYlcqf6azG0/VQZVc
tXnDsPFDHJ7gxmTeB/EA4hRL2zgOKdCzvWh2ffCMUpnhq+NyDGeVeR1zfWlGWAqk2jecnkzTIo/b
VGw7cqq10SIu88aqiQMss40QMR1Qu7tAyjmcFqe4MIckfL3xSHFizQllGL0EThbaA13LaO7jSH4w
iIqLd7DUmTU+WTAw2gb61QtVbrIlqpYvpkH5/zMhh92kKzgizrOslPsFB959njE2R/GaqAxPkXq1
DU9exkN35S0eI7nEv7Y7VHE9/b5OVu3ZZbekOreJpuo52n1l8sxc+4ATmTQ2Ht4PYUBh9n5/RgM3
rFQDROOuqeK3PZOOLsstQjG6oQ+9TXexhSK8Rhuxz141XIPVpkE4ankJN8sqZ4E58Hb/Sgm82Rdq
+70ZW3eveMaJ9lSQohMfdDZmbYBDnF45b+HNUSVVaZqz5nQ9KXu1PWBC7s6++dlAZSFYL0ZNHb8B
TVc/Yo5Ffh7R8No2UIB6JxIFC7XY61Eh2gYUTap6qLG1+rDcsyRXd+rxcBvGrTbEpJI4fMBPARWq
itVOqSkAwqvdrX6RRICQWu32zVxWYCmlHErYnV9bgu7dAFyYmBq9Ege5OTU2DZwEdJJYDq0AkwWm
aWjCdZHbUNhoPZnBhXjYu4qWr3fctY0yzPWza1TYegvU7sWtdQhA2rqtJdw8UaUIzgdS4z+9bAWS
+hI9LUyNX1Yu8IDay7kQ8/T0XopIGLaAnIUJCu0o929o1/8j7JmkQ3SfH3ZsXmE=
`protect end_protected
